DEPTH =  10240;
WIDTH =  15;
ADDRESS_RADIX = OCT;
DATA_RADIX = OCT;

CONTENT BEGIN

0000 : 00004;
0001 : 14054;
0002 : 14003;
0003 : 14004;
0004 : 50017;
0005 : 14006;
0006 : 14007;
0007 : 14010;
0010 : 14011;
0011 : 14012;
0012 : 14013;
0013 : 14014;
0014 : 14015;
0015 : 14016;
0016 : 14017;
0017 : 14020;
0020 : 50017;
0021 : 14022;
0022 : 14023;
0023 : 14024;
0024 : 50017;
0025 : 14026;
0026 : 14027;
0027 : 14030;
0030 : 50017;
0031 : 14032;
0032 : 14033;
0033 : 14034;
0034 : 50017;
0035 : 14036;
0036 : 14037;
0037 : 14040;
0040 : 50017;
0041 : 14042;
0042 : 14043;
0043 : 14044;
0044 : 50017;
0045 : 14046;
0046 : 14047;
0047 : 14050;
0050 : 50017;
0051 : 14052;
0052 : 14053;
0053 : 14054;
0054 : 34072;
0055 : 50000;
0056 : 04060;
0057 : 14060;
0060 : 04064;
0061 : 04064;
0062 : 04065;
0063 : 04064;
0064 : 64073;
0065 : 64071;
0066 : 00006;
0067 : 30051;
0070 : 00000;
0071 : 00001;
0072 : 00002;
0073 : 00004;
0074 : 00000;
0075 : 00000;
0076 : 00000;
0077 : 00000;
0100 : 00000;
0101 : 00000;
0102 : 00000;
0103 : 00000;
0104 : 00000;
0105 : 00000;
0106 : 00000;
0107 : 00000;
0110 : 00000;
0111 : 00000;
0112 : 00000;
0113 : 00000;
0114 : 00000;
0115 : 00000;
0116 : 00000;
0117 : 00000;
0120 : 00000;
0121 : 00000;
0122 : 00000;
0123 : 00000;
0124 : 00000;
0125 : 00000;
0126 : 00000;
0127 : 00000;
0130 : 00000;
0131 : 00000;
0132 : 00000;
0133 : 00000;
0134 : 00000;
0135 : 00000;
0136 : 00000;
0137 : 00000;
0140 : 00000;
0141 : 00000;
0142 : 00000;
0143 : 00000;
0144 : 00000;
0145 : 00000;
0146 : 00000;
0147 : 00000;
0150 : 00000;
0151 : 00000;
0152 : 00000;
0153 : 00000;
0154 : 00000;
0155 : 00000;
0156 : 00000;
0157 : 00000;
0160 : 00000;
0161 : 00000;
0162 : 00000;
0163 : 00000;
0164 : 00000;
0165 : 00000;
0166 : 00000;
0167 : 00000;
0170 : 00000;
0171 : 00000;
0172 : 00000;
0173 : 00000;
0174 : 00000;
0175 : 00000;
0176 : 00000;
0177 : 00000;
0200 : 00000;
0201 : 00000;
0202 : 00000;
0203 : 00000;
0204 : 00000;
0205 : 00000;
0206 : 00000;
0207 : 00000;
0210 : 00000;
0211 : 00000;
0212 : 00000;
0213 : 00000;
0214 : 00000;
0215 : 00000;
0216 : 00000;
0217 : 00000;
0220 : 00000;
0221 : 00000;
0222 : 00000;
0223 : 00000;
0224 : 00000;
0225 : 00000;
0226 : 00000;
0227 : 00000;
0230 : 00000;
0231 : 00000;
0232 : 00000;
0233 : 00000;
0234 : 00000;
0235 : 00000;
0236 : 00000;
0237 : 00000;
0240 : 00000;
0241 : 00000;
0242 : 00000;
0243 : 00000;
0244 : 00000;
0245 : 00000;
0246 : 00000;
0247 : 00000;
0250 : 00000;
0251 : 00000;
0252 : 00000;
0253 : 00000;
0254 : 00000;
0255 : 00000;
0256 : 00000;
0257 : 00000;
0260 : 00000;
0261 : 00000;
0262 : 00000;
0263 : 00000;
0264 : 00000;
0265 : 00000;
0266 : 00000;
0267 : 00000;
0270 : 00000;
0271 : 00000;
0272 : 00000;
0273 : 00000;
0274 : 00000;
0275 : 00000;
0276 : 00000;
0277 : 00000;
0300 : 00000;
0301 : 00000;
0302 : 00000;
0303 : 00000;
0304 : 00000;
0305 : 00000;
0306 : 00000;
0307 : 00000;
0310 : 00000;
0311 : 00000;
0312 : 00000;
0313 : 00000;
0314 : 00000;
0315 : 00000;
0316 : 00000;
0317 : 00000;
0320 : 00000;
0321 : 00000;
0322 : 00000;
0323 : 00000;
0324 : 00000;
0325 : 00000;
0326 : 00000;
0327 : 00000;
0330 : 00000;
0331 : 00000;
0332 : 00000;
0333 : 00000;
0334 : 00000;
0335 : 00000;
0336 : 00000;
0337 : 00000;
0340 : 00000;
0341 : 00000;
0342 : 00000;
0343 : 00000;
0344 : 00000;
0345 : 00000;
0346 : 00000;
0347 : 00000;
0350 : 00000;
0351 : 00000;
0352 : 00000;
0353 : 00000;
0354 : 00000;
0355 : 00000;
0356 : 00000;
0357 : 00000;
0360 : 00000;
0361 : 00000;
0362 : 00000;
0363 : 00000;
0364 : 00000;
0365 : 00000;
0366 : 00000;
0367 : 00000;
0370 : 00000;
0371 : 00000;
0372 : 00000;
0373 : 00000;
0374 : 00000;
0375 : 00000;
0376 : 00000;
0377 : 00000;
0400 : 00000;
0401 : 00000;
0402 : 00000;
0403 : 00000;
0404 : 00000;
0405 : 00000;
0406 : 00000;
0407 : 00000;
0410 : 00000;
0411 : 00000;
0412 : 00000;
0413 : 00000;
0414 : 00000;
0415 : 00000;
0416 : 00000;
0417 : 00000;
0420 : 00000;
0421 : 00000;
0422 : 00000;
0423 : 00000;
0424 : 00000;
0425 : 00000;
0426 : 00000;
0427 : 00000;
0430 : 00000;
0431 : 00000;
0432 : 00000;
0433 : 00000;
0434 : 00000;
0435 : 00000;
0436 : 00000;
0437 : 00000;
0440 : 00000;
0441 : 00000;
0442 : 00000;
0443 : 00000;
0444 : 00000;
0445 : 00000;
0446 : 00000;
0447 : 00000;
0450 : 00000;
0451 : 00000;
0452 : 00000;
0453 : 00000;
0454 : 00000;
0455 : 00000;
0456 : 00000;
0457 : 00000;
0460 : 00000;
0461 : 00000;
0462 : 00000;
0463 : 00000;
0464 : 00000;
0465 : 00000;
0466 : 00000;
0467 : 00000;
0470 : 00000;
0471 : 00000;
0472 : 00000;
0473 : 00000;
0474 : 00000;
0475 : 00000;
0476 : 00000;
0477 : 00000;
0500 : 00000;
0501 : 00000;
0502 : 00000;
0503 : 00000;
0504 : 00000;
0505 : 00000;
0506 : 00000;
0507 : 00000;
0510 : 00000;
0511 : 00000;
0512 : 00000;
0513 : 00000;
0514 : 00000;
0515 : 00000;
0516 : 00000;
0517 : 00000;
0520 : 00000;
0521 : 00000;
0522 : 00000;
0523 : 00000;
0524 : 00000;
0525 : 00000;
0526 : 00000;
0527 : 00000;
0530 : 00000;
0531 : 00000;
0532 : 00000;
0533 : 00000;
0534 : 00000;
0535 : 00000;
0536 : 00000;
0537 : 00000;
0540 : 00000;
0541 : 00000;
0542 : 00000;
0543 : 00000;
0544 : 00000;
0545 : 00000;
0546 : 00000;
0547 : 00000;
0550 : 00000;
0551 : 00000;
0552 : 00000;
0553 : 00000;
0554 : 00000;
0555 : 00000;
0556 : 00000;
0557 : 00000;
0560 : 00000;
0561 : 00000;
0562 : 00000;
0563 : 00000;
0564 : 00000;
0565 : 00000;
0566 : 00000;
0567 : 00000;
0570 : 00000;
0571 : 00000;
0572 : 00000;
0573 : 00000;
0574 : 00000;
0575 : 00000;
0576 : 00000;
0577 : 00000;
0600 : 00000;
0601 : 00000;
0602 : 00000;
0603 : 00000;
0604 : 00000;
0605 : 00000;
0606 : 00000;
0607 : 00000;
0610 : 00000;
0611 : 00000;
0612 : 00000;
0613 : 00000;
0614 : 00000;
0615 : 00000;
0616 : 00000;
0617 : 00000;
0620 : 00000;
0621 : 00000;
0622 : 00000;
0623 : 00000;
0624 : 00000;
0625 : 00000;
0626 : 00000;
0627 : 00000;
0630 : 00000;
0631 : 00000;
0632 : 00000;
0633 : 00000;
0634 : 00000;
0635 : 00000;
0636 : 00000;
0637 : 00000;
0640 : 00000;
0641 : 00000;
0642 : 00000;
0643 : 00000;
0644 : 00000;
0645 : 00000;
0646 : 00000;
0647 : 00000;
0650 : 00000;
0651 : 00000;
0652 : 00000;
0653 : 00000;
0654 : 00000;
0655 : 00000;
0656 : 00000;
0657 : 00000;
0660 : 00000;
0661 : 00000;
0662 : 00000;
0663 : 00000;
0664 : 00000;
0665 : 00000;
0666 : 00000;
0667 : 00000;
0670 : 00000;
0671 : 00000;
0672 : 00000;
0673 : 00000;
0674 : 00000;
0675 : 00000;
0676 : 00000;
0677 : 00000;
0700 : 00000;
0701 : 00000;
0702 : 00000;
0703 : 00000;
0704 : 00000;
0705 : 00000;
0706 : 00000;
0707 : 00000;
0710 : 00000;
0711 : 00000;
0712 : 00000;
0713 : 00000;
0714 : 00000;
0715 : 00000;
0716 : 00000;
0717 : 00000;
0720 : 00000;
0721 : 00000;
0722 : 00000;
0723 : 00000;
0724 : 00000;
0725 : 00000;
0726 : 00000;
0727 : 00000;
0730 : 00000;
0731 : 00000;
0732 : 00000;
0733 : 00000;
0734 : 00000;
0735 : 00000;
0736 : 00000;
0737 : 00000;
0740 : 00000;
0741 : 00000;
0742 : 00000;
0743 : 00000;
0744 : 00000;
0745 : 00000;
0746 : 00000;
0747 : 00000;
0750 : 00000;
0751 : 00000;
0752 : 00000;
0753 : 00000;
0754 : 00000;
0755 : 00000;
0756 : 00000;
0757 : 00000;
0760 : 00000;
0761 : 00000;
0762 : 00000;
0763 : 00000;
0764 : 00000;
0765 : 00000;
0766 : 00000;
0767 : 00000;
0770 : 00000;
0771 : 00000;
0772 : 00000;
0773 : 00000;
0774 : 00000;
0775 : 00000;
0776 : 00000;
0777 : 00000;
1000 : 00000;
1001 : 00000;
1002 : 00000;
1003 : 00000;
1004 : 00000;
1005 : 00000;
1006 : 00000;
1007 : 00000;
1010 : 00000;
1011 : 00000;
1012 : 00000;
1013 : 00000;
1014 : 00000;
1015 : 00000;
1016 : 00000;
1017 : 00000;
1020 : 00000;
1021 : 00000;
1022 : 00000;
1023 : 00000;
1024 : 00000;
1025 : 00000;
1026 : 00000;
1027 : 00000;
1030 : 00000;
1031 : 00000;
1032 : 00000;
1033 : 00000;
1034 : 00000;
1035 : 00000;
1036 : 00000;
1037 : 00000;
1040 : 00000;
1041 : 00000;
1042 : 00000;
1043 : 00000;
1044 : 00000;
1045 : 00000;
1046 : 00000;
1047 : 00000;
1050 : 00000;
1051 : 00000;
1052 : 00000;
1053 : 00000;
1054 : 00000;
1055 : 00000;
1056 : 00000;
1057 : 00000;
1060 : 00000;
1061 : 00000;
1062 : 00000;
1063 : 00000;
1064 : 00000;
1065 : 00000;
1066 : 00000;
1067 : 00000;
1070 : 00000;
1071 : 00000;
1072 : 00000;
1073 : 00000;
1074 : 00000;
1075 : 00000;
1076 : 00000;
1077 : 00000;
1100 : 00000;
1101 : 00000;
1102 : 00000;
1103 : 00000;
1104 : 00000;
1105 : 00000;
1106 : 00000;
1107 : 00000;
1110 : 00000;
1111 : 00000;
1112 : 00000;
1113 : 00000;
1114 : 00000;
1115 : 00000;
1116 : 00000;
1117 : 00000;
1120 : 00000;
1121 : 00000;
1122 : 00000;
1123 : 00000;
1124 : 00000;
1125 : 00000;
1126 : 00000;
1127 : 00000;
1130 : 00000;
1131 : 00000;
1132 : 00000;
1133 : 00000;
1134 : 00000;
1135 : 00000;
1136 : 00000;
1137 : 00000;
1140 : 00000;
1141 : 00000;
1142 : 00000;
1143 : 00000;
1144 : 00000;
1145 : 00000;
1146 : 00000;
1147 : 00000;
1150 : 00000;
1151 : 00000;
1152 : 00000;
1153 : 00000;
1154 : 00000;
1155 : 00000;
1156 : 00000;
1157 : 00000;
1160 : 00000;
1161 : 00000;
1162 : 00000;
1163 : 00000;
1164 : 00000;
1165 : 00000;
1166 : 00000;
1167 : 00000;
1170 : 00000;
1171 : 00000;
1172 : 00000;
1173 : 00000;
1174 : 00000;
1175 : 00000;
1176 : 00000;
1177 : 00000;
1200 : 00000;
1201 : 00000;
1202 : 00000;
1203 : 00000;
1204 : 00000;
1205 : 00000;
1206 : 00000;
1207 : 00000;
1210 : 00000;
1211 : 00000;
1212 : 00000;
1213 : 00000;
1214 : 00000;
1215 : 00000;
1216 : 00000;
1217 : 00000;
1220 : 00000;
1221 : 00000;
1222 : 00000;
1223 : 00000;
1224 : 00000;
1225 : 00000;
1226 : 00000;
1227 : 00000;
1230 : 00000;
1231 : 00000;
1232 : 00000;
1233 : 00000;
1234 : 00000;
1235 : 00000;
1236 : 00000;
1237 : 00000;
1240 : 00000;
1241 : 00000;
1242 : 00000;
1243 : 00000;
1244 : 00000;
1245 : 00000;
1246 : 00000;
1247 : 00000;
1250 : 00000;
1251 : 00000;
1252 : 00000;
1253 : 00000;
1254 : 00000;
1255 : 00000;
1256 : 00000;
1257 : 00000;
1260 : 00000;
1261 : 00000;
1262 : 00000;
1263 : 00000;
1264 : 00000;
1265 : 00000;
1266 : 00000;
1267 : 00000;
1270 : 00000;
1271 : 00000;
1272 : 00000;
1273 : 00000;
1274 : 00000;
1275 : 00000;
1276 : 00000;
1277 : 00000;
1300 : 00000;
1301 : 00000;
1302 : 00000;
1303 : 00000;
1304 : 00000;
1305 : 00000;
1306 : 00000;
1307 : 00000;
1310 : 00000;
1311 : 00000;
1312 : 00000;
1313 : 00000;
1314 : 00000;
1315 : 00000;
1316 : 00000;
1317 : 00000;
1320 : 00000;
1321 : 00000;
1322 : 00000;
1323 : 00000;
1324 : 00000;
1325 : 00000;
1326 : 00000;
1327 : 00000;
1330 : 00000;
1331 : 00000;
1332 : 00000;
1333 : 00000;
1334 : 00000;
1335 : 00000;
1336 : 00000;
1337 : 00000;
1340 : 00000;
1341 : 00000;
1342 : 00000;
1343 : 00000;
1344 : 00000;
1345 : 00000;
1346 : 00000;
1347 : 00000;
1350 : 00000;
1351 : 00000;
1352 : 00000;
1353 : 00000;
1354 : 00000;
1355 : 00000;
1356 : 00000;
1357 : 00000;
1360 : 00000;
1361 : 00000;
1362 : 00000;
1363 : 00000;
1364 : 00000;
1365 : 00000;
1366 : 00000;
1367 : 00000;
1370 : 00000;
1371 : 00000;
1372 : 00000;
1373 : 00000;
1374 : 00000;
1375 : 00000;
1376 : 00000;
1377 : 00000;
1400 : 00000;
1401 : 00000;
1402 : 00000;
1403 : 00000;
1404 : 00000;
1405 : 00000;
1406 : 00000;
1407 : 00000;
1410 : 00000;
1411 : 00000;
1412 : 00000;
1413 : 00000;
1414 : 00000;
1415 : 00000;
1416 : 00000;
1417 : 00000;
1420 : 00000;
1421 : 00000;
1422 : 00000;
1423 : 00000;
1424 : 00000;
1425 : 00000;
1426 : 00000;
1427 : 00000;
1430 : 00000;
1431 : 00000;
1432 : 00000;
1433 : 00000;
1434 : 00000;
1435 : 00000;
1436 : 00000;
1437 : 00000;
1440 : 00000;
1441 : 00000;
1442 : 00000;
1443 : 00000;
1444 : 00000;
1445 : 00000;
1446 : 00000;
1447 : 00000;
1450 : 00000;
1451 : 00000;
1452 : 00000;
1453 : 00000;
1454 : 00000;
1455 : 00000;
1456 : 00000;
1457 : 00000;
1460 : 00000;
1461 : 00000;
1462 : 00000;
1463 : 00000;
1464 : 00000;
1465 : 00000;
1466 : 00000;
1467 : 00000;
1470 : 00000;
1471 : 00000;
1472 : 00000;
1473 : 00000;
1474 : 00000;
1475 : 00000;
1476 : 00000;
1477 : 00000;
1500 : 00000;
1501 : 00000;
1502 : 00000;
1503 : 00000;
1504 : 00000;
1505 : 00000;
1506 : 00000;
1507 : 00000;
1510 : 00000;
1511 : 00000;
1512 : 00000;
1513 : 00000;
1514 : 00000;
1515 : 00000;
1516 : 00000;
1517 : 00000;
1520 : 00000;
1521 : 00000;
1522 : 00000;
1523 : 00000;
1524 : 00000;
1525 : 00000;
1526 : 00000;
1527 : 00000;
1530 : 00000;
1531 : 00000;
1532 : 00000;
1533 : 00000;
1534 : 00000;
1535 : 00000;
1536 : 00000;
1537 : 00000;
1540 : 00000;
1541 : 00000;
1542 : 00000;
1543 : 00000;
1544 : 00000;
1545 : 00000;
1546 : 00000;
1547 : 00000;
1550 : 00000;
1551 : 00000;
1552 : 00000;
1553 : 00000;
1554 : 00000;
1555 : 00000;
1556 : 00000;
1557 : 00000;
1560 : 00000;
1561 : 00000;
1562 : 00000;
1563 : 00000;
1564 : 00000;
1565 : 00000;
1566 : 00000;
1567 : 00000;
1570 : 00000;
1571 : 00000;
1572 : 00000;
1573 : 00000;
1574 : 00000;
1575 : 00000;
1576 : 00000;
1577 : 00000;
1600 : 00000;
1601 : 00000;
1602 : 00000;
1603 : 00000;
1604 : 00000;
1605 : 00000;
1606 : 00000;
1607 : 00000;
1610 : 00000;
1611 : 00000;
1612 : 00000;
1613 : 00000;
1614 : 00000;
1615 : 00000;
1616 : 00000;
1617 : 00000;
1620 : 00000;
1621 : 00000;
1622 : 00000;
1623 : 00000;
1624 : 00000;
1625 : 00000;
1626 : 00000;
1627 : 00000;
1630 : 00000;
1631 : 00000;
1632 : 00000;
1633 : 00000;
1634 : 00000;
1635 : 00000;
1636 : 00000;
1637 : 00000;
1640 : 00000;
1641 : 00000;
1642 : 00000;
1643 : 00000;
1644 : 00000;
1645 : 00000;
1646 : 00000;
1647 : 00000;
1650 : 00000;
1651 : 00000;
1652 : 00000;
1653 : 00000;
1654 : 00000;
1655 : 00000;
1656 : 00000;
1657 : 00000;
1660 : 00000;
1661 : 00000;
1662 : 00000;
1663 : 00000;
1664 : 00000;
1665 : 00000;
1666 : 00000;
1667 : 00000;
1670 : 00000;
1671 : 00000;
1672 : 00000;
1673 : 00000;
1674 : 00000;
1675 : 00000;
1676 : 00000;
1677 : 00000;
1700 : 00000;
1701 : 00000;
1702 : 00000;
1703 : 00000;
1704 : 00000;
1705 : 00000;
1706 : 00000;
1707 : 00000;
1710 : 00000;
1711 : 00000;
1712 : 00000;
1713 : 00000;
1714 : 00000;
1715 : 00000;
1716 : 00000;
1717 : 00000;
1720 : 00000;
1721 : 00000;
1722 : 00000;
1723 : 00000;
1724 : 00000;
1725 : 00000;
1726 : 00000;
1727 : 00000;
1730 : 00000;
1731 : 00000;
1732 : 00000;
1733 : 00000;
1734 : 00000;
1735 : 00000;
1736 : 00000;
1737 : 00000;
1740 : 00000;
1741 : 00000;
1742 : 00000;
1743 : 00000;
1744 : 00000;
1745 : 00000;
1746 : 00000;
1747 : 00000;
1750 : 00000;
1751 : 00000;
1752 : 00000;
1753 : 00000;
1754 : 00000;
1755 : 00000;
1756 : 00000;
1757 : 00000;
1760 : 00000;
1761 : 00000;
1762 : 00000;
1763 : 00000;
1764 : 00000;
1765 : 00000;
1766 : 00000;
1767 : 00000;
1770 : 00000;
1771 : 00000;
1772 : 00000;
1773 : 00000;
1774 : 00000;
1775 : 00000;
1776 : 00000;
1777 : 00000;
2000 : 00000;
2001 : 00000;
2002 : 00000;
2003 : 00000;
2004 : 00000;
2005 : 00000;
2006 : 00000;
2007 : 00000;
2010 : 00000;
2011 : 00000;
2012 : 00000;
2013 : 00000;
2014 : 00000;
2015 : 00000;
2016 : 00000;
2017 : 00000;
2020 : 00000;
2021 : 00000;
2022 : 00000;
2023 : 00000;
2024 : 00000;
2025 : 00000;
2026 : 00000;
2027 : 00000;
2030 : 00000;
2031 : 00000;
2032 : 00000;
2033 : 00000;
2034 : 00000;
2035 : 00000;
2036 : 00000;
2037 : 00000;
2040 : 00000;
2041 : 00000;
2042 : 00000;
2043 : 00000;
2044 : 00000;
2045 : 00000;
2046 : 00000;
2047 : 00000;
2050 : 00000;
2051 : 00000;
2052 : 00000;
2053 : 00000;
2054 : 00000;
2055 : 00000;
2056 : 00000;
2057 : 00000;
2060 : 00000;
2061 : 00000;
2062 : 00000;
2063 : 00000;
2064 : 00000;
2065 : 00000;
2066 : 00000;
2067 : 00000;
2070 : 00000;
2071 : 00000;
2072 : 00000;
2073 : 00000;
2074 : 00000;
2075 : 00000;
2076 : 00000;
2077 : 00000;
2100 : 00000;
2101 : 00000;
2102 : 00000;
2103 : 00000;
2104 : 00000;
2105 : 00000;
2106 : 00000;
2107 : 00000;
2110 : 00000;
2111 : 00000;
2112 : 00000;
2113 : 00000;
2114 : 00000;
2115 : 00000;
2116 : 00000;
2117 : 00000;
2120 : 00000;
2121 : 00000;
2122 : 00000;
2123 : 00000;
2124 : 00000;
2125 : 00000;
2126 : 00000;
2127 : 00000;
2130 : 00000;
2131 : 00000;
2132 : 00000;
2133 : 00000;
2134 : 00000;
2135 : 00000;
2136 : 00000;
2137 : 00000;
2140 : 00000;
2141 : 00000;
2142 : 00000;
2143 : 00000;
2144 : 00000;
2145 : 00000;
2146 : 00000;
2147 : 00000;
2150 : 00000;
2151 : 00000;
2152 : 00000;
2153 : 00000;
2154 : 00000;
2155 : 00000;
2156 : 00000;
2157 : 00000;
2160 : 00000;
2161 : 00000;
2162 : 00000;
2163 : 00000;
2164 : 00000;
2165 : 00000;
2166 : 00000;
2167 : 00000;
2170 : 00000;
2171 : 00000;
2172 : 00000;
2173 : 00000;
2174 : 00000;
2175 : 00000;
2176 : 00000;
2177 : 00000;
2200 : 00000;
2201 : 00000;
2202 : 00000;
2203 : 00000;
2204 : 00000;
2205 : 00000;
2206 : 00000;
2207 : 00000;
2210 : 00000;
2211 : 00000;
2212 : 00000;
2213 : 00000;
2214 : 00000;
2215 : 00000;
2216 : 00000;
2217 : 00000;
2220 : 00000;
2221 : 00000;
2222 : 00000;
2223 : 00000;
2224 : 00000;
2225 : 00000;
2226 : 00000;
2227 : 00000;
2230 : 00000;
2231 : 00000;
2232 : 00000;
2233 : 00000;
2234 : 00000;
2235 : 00000;
2236 : 00000;
2237 : 00000;
2240 : 00000;
2241 : 00000;
2242 : 00000;
2243 : 00000;
2244 : 00000;
2245 : 00000;
2246 : 00000;
2247 : 00000;
2250 : 00000;
2251 : 00000;
2252 : 00000;
2253 : 00000;
2254 : 00000;
2255 : 00000;
2256 : 00000;
2257 : 00000;
2260 : 00000;
2261 : 00000;
2262 : 00000;
2263 : 00000;
2264 : 00000;
2265 : 00000;
2266 : 00000;
2267 : 00000;
2270 : 00000;
2271 : 00000;
2272 : 00000;
2273 : 00000;
2274 : 00000;
2275 : 00000;
2276 : 00000;
2277 : 00000;
2300 : 00000;
2301 : 00000;
2302 : 00000;
2303 : 00000;
2304 : 00000;
2305 : 00000;
2306 : 00000;
2307 : 00000;
2310 : 00000;
2311 : 00000;
2312 : 00000;
2313 : 00000;
2314 : 00000;
2315 : 00000;
2316 : 00000;
2317 : 00000;
2320 : 00000;
2321 : 00000;
2322 : 00000;
2323 : 00000;
2324 : 00000;
2325 : 00000;
2326 : 00000;
2327 : 00000;
2330 : 00000;
2331 : 00000;
2332 : 00000;
2333 : 00000;
2334 : 00000;
2335 : 00000;
2336 : 00000;
2337 : 00000;
2340 : 00000;
2341 : 00000;
2342 : 00000;
2343 : 00000;
2344 : 00000;
2345 : 00000;
2346 : 00000;
2347 : 00000;
2350 : 00000;
2351 : 00000;
2352 : 00000;
2353 : 00000;
2354 : 00000;
2355 : 00000;
2356 : 00000;
2357 : 00000;
2360 : 00000;
2361 : 00000;
2362 : 00000;
2363 : 00000;
2364 : 00000;
2365 : 00000;
2366 : 00000;
2367 : 00000;
2370 : 00000;
2371 : 00000;
2372 : 00000;
2373 : 00000;
2374 : 00000;
2375 : 00000;
2376 : 00000;
2377 : 00000;
2400 : 00000;
2401 : 00000;
2402 : 00000;
2403 : 00000;
2404 : 00000;
2405 : 00000;
2406 : 00000;
2407 : 00000;
2410 : 00000;
2411 : 00000;
2412 : 00000;
2413 : 00000;
2414 : 00000;
2415 : 00000;
2416 : 00000;
2417 : 00000;
2420 : 00000;
2421 : 00000;
2422 : 00000;
2423 : 00000;
2424 : 00000;
2425 : 00000;
2426 : 00000;
2427 : 00000;
2430 : 00000;
2431 : 00000;
2432 : 00000;
2433 : 00000;
2434 : 00000;
2435 : 00000;
2436 : 00000;
2437 : 00000;
2440 : 00000;
2441 : 00000;
2442 : 00000;
2443 : 00000;
2444 : 00000;
2445 : 00000;
2446 : 00000;
2447 : 00000;
2450 : 00000;
2451 : 00000;
2452 : 00000;
2453 : 00000;
2454 : 00000;
2455 : 00000;
2456 : 00000;
2457 : 00000;
2460 : 00000;
2461 : 00000;
2462 : 00000;
2463 : 00000;
2464 : 00000;
2465 : 00000;
2466 : 00000;
2467 : 00000;
2470 : 00000;
2471 : 00000;
2472 : 00000;
2473 : 00000;
2474 : 00000;
2475 : 00000;
2476 : 00000;
2477 : 00000;
2500 : 00000;
2501 : 00000;
2502 : 00000;
2503 : 00000;
2504 : 00000;
2505 : 00000;
2506 : 00000;
2507 : 00000;
2510 : 00000;
2511 : 00000;
2512 : 00000;
2513 : 00000;
2514 : 00000;
2515 : 00000;
2516 : 00000;
2517 : 00000;
2520 : 00000;
2521 : 00000;
2522 : 00000;
2523 : 00000;
2524 : 00000;
2525 : 00000;
2526 : 00000;
2527 : 00000;
2530 : 00000;
2531 : 00000;
2532 : 00000;
2533 : 00000;
2534 : 00000;
2535 : 00000;
2536 : 00000;
2537 : 00000;
2540 : 00000;
2541 : 00000;
2542 : 00000;
2543 : 00000;
2544 : 00000;
2545 : 00000;
2546 : 00000;
2547 : 00000;
2550 : 00000;
2551 : 00000;
2552 : 00000;
2553 : 00000;
2554 : 00000;
2555 : 00000;
2556 : 00000;
2557 : 00000;
2560 : 00000;
2561 : 00000;
2562 : 00000;
2563 : 00000;
2564 : 00000;
2565 : 00000;
2566 : 00000;
2567 : 00000;
2570 : 00000;
2571 : 00000;
2572 : 00000;
2573 : 00000;
2574 : 00000;
2575 : 00000;
2576 : 00000;
2577 : 00000;
2600 : 00000;
2601 : 00000;
2602 : 00000;
2603 : 00000;
2604 : 00000;
2605 : 00000;
2606 : 00000;
2607 : 00000;
2610 : 00000;
2611 : 00000;
2612 : 00000;
2613 : 00000;
2614 : 00000;
2615 : 00000;
2616 : 00000;
2617 : 00000;
2620 : 00000;
2621 : 00000;
2622 : 00000;
2623 : 00000;
2624 : 00000;
2625 : 00000;
2626 : 00000;
2627 : 00000;
2630 : 00000;
2631 : 00000;
2632 : 00000;
2633 : 00000;
2634 : 00000;
2635 : 00000;
2636 : 00000;
2637 : 00000;
2640 : 00000;
2641 : 00000;
2642 : 00000;
2643 : 00000;
2644 : 00000;
2645 : 00000;
2646 : 00000;
2647 : 00000;
2650 : 00000;
2651 : 00000;
2652 : 00000;
2653 : 00000;
2654 : 00000;
2655 : 00000;
2656 : 00000;
2657 : 00000;
2660 : 00000;
2661 : 00000;
2662 : 00000;
2663 : 00000;
2664 : 00000;
2665 : 00000;
2666 : 00000;
2667 : 00000;
2670 : 00000;
2671 : 00000;
2672 : 00000;
2673 : 00000;
2674 : 00000;
2675 : 00000;
2676 : 00000;
2677 : 00000;
2700 : 00000;
2701 : 00000;
2702 : 00000;
2703 : 00000;
2704 : 00000;
2705 : 00000;
2706 : 00000;
2707 : 00000;
2710 : 00000;
2711 : 00000;
2712 : 00000;
2713 : 00000;
2714 : 00000;
2715 : 00000;
2716 : 00000;
2717 : 00000;
2720 : 00000;
2721 : 00000;
2722 : 00000;
2723 : 00000;
2724 : 00000;
2725 : 00000;
2726 : 00000;
2727 : 00000;
2730 : 00000;
2731 : 00000;
2732 : 00000;
2733 : 00000;
2734 : 00000;
2735 : 00000;
2736 : 00000;
2737 : 00000;
2740 : 00000;
2741 : 00000;
2742 : 00000;
2743 : 00000;
2744 : 00000;
2745 : 00000;
2746 : 00000;
2747 : 00000;
2750 : 00000;
2751 : 00000;
2752 : 00000;
2753 : 00000;
2754 : 00000;
2755 : 00000;
2756 : 00000;
2757 : 00000;
2760 : 00000;
2761 : 00000;
2762 : 00000;
2763 : 00000;
2764 : 00000;
2765 : 00000;
2766 : 00000;
2767 : 00000;
2770 : 00000;
2771 : 00000;
2772 : 00000;
2773 : 00000;
2774 : 00000;
2775 : 00000;
2776 : 00000;
2777 : 00000;
3000 : 00000;
3001 : 00000;
3002 : 00000;
3003 : 00000;
3004 : 00000;
3005 : 00000;
3006 : 00000;
3007 : 00000;
3010 : 00000;
3011 : 00000;
3012 : 00000;
3013 : 00000;
3014 : 00000;
3015 : 00000;
3016 : 00000;
3017 : 00000;
3020 : 00000;
3021 : 00000;
3022 : 00000;
3023 : 00000;
3024 : 00000;
3025 : 00000;
3026 : 00000;
3027 : 00000;
3030 : 00000;
3031 : 00000;
3032 : 00000;
3033 : 00000;
3034 : 00000;
3035 : 00000;
3036 : 00000;
3037 : 00000;
3040 : 00000;
3041 : 00000;
3042 : 00000;
3043 : 00000;
3044 : 00000;
3045 : 00000;
3046 : 00000;
3047 : 00000;
3050 : 00000;
3051 : 00000;
3052 : 00000;
3053 : 00000;
3054 : 00000;
3055 : 00000;
3056 : 00000;
3057 : 00000;
3060 : 00000;
3061 : 00000;
3062 : 00000;
3063 : 00000;
3064 : 00000;
3065 : 00000;
3066 : 00000;
3067 : 00000;
3070 : 00000;
3071 : 00000;
3072 : 00000;
3073 : 00000;
3074 : 00000;
3075 : 00000;
3076 : 00000;
3077 : 00000;
3100 : 00000;
3101 : 00000;
3102 : 00000;
3103 : 00000;
3104 : 00000;
3105 : 00000;
3106 : 00000;
3107 : 00000;
3110 : 00000;
3111 : 00000;
3112 : 00000;
3113 : 00000;
3114 : 00000;
3115 : 00000;
3116 : 00000;
3117 : 00000;
3120 : 00000;
3121 : 00000;
3122 : 00000;
3123 : 00000;
3124 : 00000;
3125 : 00000;
3126 : 00000;
3127 : 00000;
3130 : 00000;
3131 : 00000;
3132 : 00000;
3133 : 00000;
3134 : 00000;
3135 : 00000;
3136 : 00000;
3137 : 00000;
3140 : 00000;
3141 : 00000;
3142 : 00000;
3143 : 00000;
3144 : 00000;
3145 : 00000;
3146 : 00000;
3147 : 00000;
3150 : 00000;
3151 : 00000;
3152 : 00000;
3153 : 00000;
3154 : 00000;
3155 : 00000;
3156 : 00000;
3157 : 00000;
3160 : 00000;
3161 : 00000;
3162 : 00000;
3163 : 00000;
3164 : 00000;
3165 : 00000;
3166 : 00000;
3167 : 00000;
3170 : 00000;
3171 : 00000;
3172 : 00000;
3173 : 00000;
3174 : 00000;
3175 : 00000;
3176 : 00000;
3177 : 00000;
3200 : 00000;
3201 : 00000;
3202 : 00000;
3203 : 00000;
3204 : 00000;
3205 : 00000;
3206 : 00000;
3207 : 00000;
3210 : 00000;
3211 : 00000;
3212 : 00000;
3213 : 00000;
3214 : 00000;
3215 : 00000;
3216 : 00000;
3217 : 00000;
3220 : 00000;
3221 : 00000;
3222 : 00000;
3223 : 00000;
3224 : 00000;
3225 : 00000;
3226 : 00000;
3227 : 00000;
3230 : 00000;
3231 : 00000;
3232 : 00000;
3233 : 00000;
3234 : 00000;
3235 : 00000;
3236 : 00000;
3237 : 00000;
3240 : 00000;
3241 : 00000;
3242 : 00000;
3243 : 00000;
3244 : 00000;
3245 : 00000;
3246 : 00000;
3247 : 00000;
3250 : 00000;
3251 : 00000;
3252 : 00000;
3253 : 00000;
3254 : 00000;
3255 : 00000;
3256 : 00000;
3257 : 00000;
3260 : 00000;
3261 : 00000;
3262 : 00000;
3263 : 00000;
3264 : 00000;
3265 : 00000;
3266 : 00000;
3267 : 00000;
3270 : 00000;
3271 : 00000;
3272 : 00000;
3273 : 00000;
3274 : 00000;
3275 : 00000;
3276 : 00000;
3277 : 00000;
3300 : 00000;
3301 : 00000;
3302 : 00000;
3303 : 00000;
3304 : 00000;
3305 : 00000;
3306 : 00000;
3307 : 00000;
3310 : 00000;
3311 : 00000;
3312 : 00000;
3313 : 00000;
3314 : 00000;
3315 : 00000;
3316 : 00000;
3317 : 00000;
3320 : 00000;
3321 : 00000;
3322 : 00000;
3323 : 00000;
3324 : 00000;
3325 : 00000;
3326 : 00000;
3327 : 00000;
3330 : 00000;
3331 : 00000;
3332 : 00000;
3333 : 00000;
3334 : 00000;
3335 : 00000;
3336 : 00000;
3337 : 00000;
3340 : 00000;
3341 : 00000;
3342 : 00000;
3343 : 00000;
3344 : 00000;
3345 : 00000;
3346 : 00000;
3347 : 00000;
3350 : 00000;
3351 : 00000;
3352 : 00000;
3353 : 00000;
3354 : 00000;
3355 : 00000;
3356 : 00000;
3357 : 00000;
3360 : 00000;
3361 : 00000;
3362 : 00000;
3363 : 00000;
3364 : 00000;
3365 : 00000;
3366 : 00000;
3367 : 00000;
3370 : 00000;
3371 : 00000;
3372 : 00000;
3373 : 00000;
3374 : 00000;
3375 : 00000;
3376 : 00000;
3377 : 00000;
3400 : 00000;
3401 : 00000;
3402 : 00000;
3403 : 00000;
3404 : 00000;
3405 : 00000;
3406 : 00000;
3407 : 00000;
3410 : 00000;
3411 : 00000;
3412 : 00000;
3413 : 00000;
3414 : 00000;
3415 : 00000;
3416 : 00000;
3417 : 00000;
3420 : 00000;
3421 : 00000;
3422 : 00000;
3423 : 00000;
3424 : 00000;
3425 : 00000;
3426 : 00000;
3427 : 00000;
3430 : 00000;
3431 : 00000;
3432 : 00000;
3433 : 00000;
3434 : 00000;
3435 : 00000;
3436 : 00000;
3437 : 00000;
3440 : 00000;
3441 : 00000;
3442 : 00000;
3443 : 00000;
3444 : 00000;
3445 : 00000;
3446 : 00000;
3447 : 00000;
3450 : 00000;
3451 : 00000;
3452 : 00000;
3453 : 00000;
3454 : 00000;
3455 : 00000;
3456 : 00000;
3457 : 00000;
3460 : 00000;
3461 : 00000;
3462 : 00000;
3463 : 00000;
3464 : 00000;
3465 : 00000;
3466 : 00000;
3467 : 00000;
3470 : 00000;
3471 : 00000;
3472 : 00000;
3473 : 00000;
3474 : 00000;
3475 : 00000;
3476 : 00000;
3477 : 00000;
3500 : 00000;
3501 : 00000;
3502 : 00000;
3503 : 00000;
3504 : 00000;
3505 : 00000;
3506 : 00000;
3507 : 00000;
3510 : 00000;
3511 : 00000;
3512 : 00000;
3513 : 00000;
3514 : 00000;
3515 : 00000;
3516 : 00000;
3517 : 00000;
3520 : 00000;
3521 : 00000;
3522 : 00000;
3523 : 00000;
3524 : 00000;
3525 : 00000;
3526 : 00000;
3527 : 00000;
3530 : 00000;
3531 : 00000;
3532 : 00000;
3533 : 00000;
3534 : 00000;
3535 : 00000;
3536 : 00000;
3537 : 00000;
3540 : 00000;
3541 : 00000;
3542 : 00000;
3543 : 00000;
3544 : 00000;
3545 : 00000;
3546 : 00000;
3547 : 00000;
3550 : 00000;
3551 : 00000;
3552 : 00000;
3553 : 00000;
3554 : 00000;
3555 : 00000;
3556 : 00000;
3557 : 00000;
3560 : 00000;
3561 : 00000;
3562 : 00000;
3563 : 00000;
3564 : 00000;
3565 : 00000;
3566 : 00000;
3567 : 00000;
3570 : 00000;
3571 : 00000;
3572 : 00000;
3573 : 00000;
3574 : 00000;
3575 : 00000;
3576 : 00000;
3577 : 00000;
3600 : 00000;
3601 : 00000;
3602 : 00000;
3603 : 00000;
3604 : 00000;
3605 : 00000;
3606 : 00000;
3607 : 00000;
3610 : 00000;
3611 : 00000;
3612 : 00000;
3613 : 00000;
3614 : 00000;
3615 : 00000;
3616 : 00000;
3617 : 00000;
3620 : 00000;
3621 : 00000;
3622 : 00000;
3623 : 00000;
3624 : 00000;
3625 : 00000;
3626 : 00000;
3627 : 00000;
3630 : 00000;
3631 : 00000;
3632 : 00000;
3633 : 00000;
3634 : 00000;
3635 : 00000;
3636 : 00000;
3637 : 00000;
3640 : 00000;
3641 : 00000;
3642 : 00000;
3643 : 00000;
3644 : 00000;
3645 : 00000;
3646 : 00000;
3647 : 00000;
3650 : 00000;
3651 : 00000;
3652 : 00000;
3653 : 00000;
3654 : 00000;
3655 : 00000;
3656 : 00000;
3657 : 00000;
3660 : 00000;
3661 : 00000;
3662 : 00000;
3663 : 00000;
3664 : 00000;
3665 : 00000;
3666 : 00000;
3667 : 00000;
3670 : 00000;
3671 : 00000;
3672 : 00000;
3673 : 00000;
3674 : 00000;
3675 : 00000;
3676 : 00000;
3677 : 00000;
3700 : 00000;
3701 : 00000;
3702 : 00000;
3703 : 00000;
3704 : 00000;
3705 : 00000;
3706 : 00000;
3707 : 00000;
3710 : 00000;
3711 : 00000;
3712 : 00000;
3713 : 00000;
3714 : 00000;
3715 : 00000;
3716 : 00000;
3717 : 00000;
3720 : 00000;
3721 : 00000;
3722 : 00000;
3723 : 00000;
3724 : 00000;
3725 : 00000;
3726 : 00000;
3727 : 00000;
3730 : 00000;
3731 : 00000;
3732 : 00000;
3733 : 00000;
3734 : 00000;
3735 : 00000;
3736 : 00000;
3737 : 00000;
3740 : 00000;
3741 : 00000;
3742 : 00000;
3743 : 00000;
3744 : 00000;
3745 : 00000;
3746 : 00000;
3747 : 00000;
3750 : 00000;
3751 : 00000;
3752 : 00000;
3753 : 00000;
3754 : 00000;
3755 : 00000;
3756 : 00000;
3757 : 00000;
3760 : 00000;
3761 : 00000;
3762 : 00000;
3763 : 00000;
3764 : 00000;
3765 : 00000;
3766 : 00000;
3767 : 00000;
3770 : 00000;
3771 : 00000;
3772 : 00000;
3773 : 00000;
3774 : 00000;
3775 : 00000;
3776 : 00000;
3777 : 00000;
4000 : 00000;
4001 : 00000;
4002 : 00000;
4003 : 00000;
4004 : 00000;
4005 : 00000;
4006 : 00000;
4007 : 00000;
4010 : 00000;
4011 : 00000;
4012 : 00000;
4013 : 00000;
4014 : 00000;
4015 : 00000;
4016 : 00000;
4017 : 00000;
4020 : 00000;
4021 : 00000;
4022 : 00000;
4023 : 00000;
4024 : 00000;
4025 : 00000;
4026 : 00000;
4027 : 00000;
4030 : 00000;
4031 : 00000;
4032 : 00000;
4033 : 00000;
4034 : 00000;
4035 : 00000;
4036 : 00000;
4037 : 00000;
4040 : 00000;
4041 : 00000;
4042 : 00000;
4043 : 00000;
4044 : 00000;
4045 : 00000;
4046 : 00000;
4047 : 00000;
4050 : 00000;
4051 : 00000;
4052 : 00000;
4053 : 00000;
4054 : 00000;
4055 : 00000;
4056 : 00000;
4057 : 00000;
4060 : 00000;
4061 : 00000;
4062 : 00000;
4063 : 00000;
4064 : 00000;
4065 : 00000;
4066 : 00000;
4067 : 00000;
4070 : 00000;
4071 : 00000;
4072 : 00000;
4073 : 00000;
4074 : 00000;
4075 : 00000;
4076 : 00000;
4077 : 00000;
4100 : 00000;
4101 : 00000;
4102 : 00000;
4103 : 00000;
4104 : 00000;
4105 : 00000;
4106 : 00000;
4107 : 00000;
4110 : 00000;
4111 : 00000;
4112 : 00000;
4113 : 00000;
4114 : 00000;
4115 : 00000;
4116 : 00000;
4117 : 00000;
4120 : 00000;
4121 : 00000;
4122 : 00000;
4123 : 00000;
4124 : 00000;
4125 : 00000;
4126 : 00000;
4127 : 00000;
4130 : 00000;
4131 : 00000;
4132 : 00000;
4133 : 00000;
4134 : 00000;
4135 : 00000;
4136 : 00000;
4137 : 00000;
4140 : 00000;
4141 : 00000;
4142 : 00000;
4143 : 00000;
4144 : 00000;
4145 : 00000;
4146 : 00000;
4147 : 00000;
4150 : 00000;
4151 : 00000;
4152 : 00000;
4153 : 00000;
4154 : 00000;
4155 : 00000;
4156 : 00000;
4157 : 00000;
4160 : 00000;
4161 : 00000;
4162 : 00000;
4163 : 00000;
4164 : 00000;
4165 : 00000;
4166 : 00000;
4167 : 00000;
4170 : 00000;
4171 : 00000;
4172 : 00000;
4173 : 00000;
4174 : 00000;
4175 : 00000;
4176 : 00000;
4177 : 00000;
4200 : 00000;
4201 : 00000;
4202 : 00000;
4203 : 00000;
4204 : 00000;
4205 : 00000;
4206 : 00000;
4207 : 00000;
4210 : 00000;
4211 : 00000;
4212 : 00000;
4213 : 00000;
4214 : 00000;
4215 : 00000;
4216 : 00000;
4217 : 00000;
4220 : 00000;
4221 : 00000;
4222 : 00000;
4223 : 00000;
4224 : 00000;
4225 : 00000;
4226 : 00000;
4227 : 00000;
4230 : 00000;
4231 : 00000;
4232 : 00000;
4233 : 00000;
4234 : 00000;
4235 : 00000;
4236 : 00000;
4237 : 00000;
4240 : 00000;
4241 : 00000;
4242 : 00000;
4243 : 00000;
4244 : 00000;
4245 : 00000;
4246 : 00000;
4247 : 00000;
4250 : 00000;
4251 : 00000;
4252 : 00000;
4253 : 00000;
4254 : 00000;
4255 : 00000;
4256 : 00000;
4257 : 00000;
4260 : 00000;
4261 : 00000;
4262 : 00000;
4263 : 00000;
4264 : 00000;
4265 : 00000;
4266 : 00000;
4267 : 00000;
4270 : 00000;
4271 : 00000;
4272 : 00000;
4273 : 00000;
4274 : 00000;
4275 : 00000;
4276 : 00000;
4277 : 00000;
4300 : 00000;
4301 : 00000;
4302 : 00000;
4303 : 00000;
4304 : 00000;
4305 : 00000;
4306 : 00000;
4307 : 00000;
4310 : 00000;
4311 : 00000;
4312 : 00000;
4313 : 00000;
4314 : 00000;
4315 : 00000;
4316 : 00000;
4317 : 00000;
4320 : 00000;
4321 : 00000;
4322 : 00000;
4323 : 00000;
4324 : 00000;
4325 : 00000;
4326 : 00000;
4327 : 00000;
4330 : 00000;
4331 : 00000;
4332 : 00000;
4333 : 00000;
4334 : 00000;
4335 : 00000;
4336 : 00000;
4337 : 00000;
4340 : 00000;
4341 : 00000;
4342 : 00000;
4343 : 00000;
4344 : 00000;
4345 : 00000;
4346 : 00000;
4347 : 00000;
4350 : 00000;
4351 : 00000;
4352 : 00000;
4353 : 00000;
4354 : 00000;
4355 : 00000;
4356 : 00000;
4357 : 00000;
4360 : 00000;
4361 : 00000;
4362 : 00000;
4363 : 00000;
4364 : 00000;
4365 : 00000;
4366 : 00000;
4367 : 00000;
4370 : 00000;
4371 : 00000;
4372 : 00000;
4373 : 00000;
4374 : 00000;
4375 : 00000;
4376 : 00000;
4377 : 00000;
4400 : 00000;
4401 : 00000;
4402 : 00000;
4403 : 00000;
4404 : 00000;
4405 : 00000;
4406 : 00000;
4407 : 00000;
4410 : 00000;
4411 : 00000;
4412 : 00000;
4413 : 00000;
4414 : 00000;
4415 : 00000;
4416 : 00000;
4417 : 00000;
4420 : 00000;
4421 : 00000;
4422 : 00000;
4423 : 00000;
4424 : 00000;
4425 : 00000;
4426 : 00000;
4427 : 00000;
4430 : 00000;
4431 : 00000;
4432 : 00000;
4433 : 00000;
4434 : 00000;
4435 : 00000;
4436 : 00000;
4437 : 00000;
4440 : 00000;
4441 : 00000;
4442 : 00000;
4443 : 00000;
4444 : 00000;
4445 : 00000;
4446 : 00000;
4447 : 00000;
4450 : 00000;
4451 : 00000;
4452 : 00000;
4453 : 00000;
4454 : 00000;
4455 : 00000;
4456 : 00000;
4457 : 00000;
4460 : 00000;
4461 : 00000;
4462 : 00000;
4463 : 00000;
4464 : 00000;
4465 : 00000;
4466 : 00000;
4467 : 00000;
4470 : 00000;
4471 : 00000;
4472 : 00000;
4473 : 00000;
4474 : 00000;
4475 : 00000;
4476 : 00000;
4477 : 00000;
4500 : 00000;
4501 : 00000;
4502 : 00000;
4503 : 00000;
4504 : 00000;
4505 : 00000;
4506 : 00000;
4507 : 00000;
4510 : 00000;
4511 : 00000;
4512 : 00000;
4513 : 00000;
4514 : 00000;
4515 : 00000;
4516 : 00000;
4517 : 00000;
4520 : 00000;
4521 : 00000;
4522 : 00000;
4523 : 00000;
4524 : 00000;
4525 : 00000;
4526 : 00000;
4527 : 00000;
4530 : 00000;
4531 : 00000;
4532 : 00000;
4533 : 00000;
4534 : 00000;
4535 : 00000;
4536 : 00000;
4537 : 00000;
4540 : 00000;
4541 : 00000;
4542 : 00000;
4543 : 00000;
4544 : 00000;
4545 : 00000;
4546 : 00000;
4547 : 00000;
4550 : 00000;
4551 : 00000;
4552 : 00000;
4553 : 00000;
4554 : 00000;
4555 : 00000;
4556 : 00000;
4557 : 00000;
4560 : 00000;
4561 : 00000;
4562 : 00000;
4563 : 00000;
4564 : 00000;
4565 : 00000;
4566 : 00000;
4567 : 00000;
4570 : 00000;
4571 : 00000;
4572 : 00000;
4573 : 00000;
4574 : 00000;
4575 : 00000;
4576 : 00000;
4577 : 00000;
4600 : 00000;
4601 : 00000;
4602 : 00000;
4603 : 00000;
4604 : 00000;
4605 : 00000;
4606 : 00000;
4607 : 00000;
4610 : 00000;
4611 : 00000;
4612 : 00000;
4613 : 00000;
4614 : 00000;
4615 : 00000;
4616 : 00000;
4617 : 00000;
4620 : 00000;
4621 : 00000;
4622 : 00000;
4623 : 00000;
4624 : 00000;
4625 : 00000;
4626 : 00000;
4627 : 00000;
4630 : 00000;
4631 : 00000;
4632 : 00000;
4633 : 00000;
4634 : 00000;
4635 : 00000;
4636 : 00000;
4637 : 00000;
4640 : 00000;
4641 : 00000;
4642 : 00000;
4643 : 00000;
4644 : 00000;
4645 : 00000;
4646 : 00000;
4647 : 00000;
4650 : 00000;
4651 : 00000;
4652 : 00000;
4653 : 00000;
4654 : 00000;
4655 : 00000;
4656 : 00000;
4657 : 00000;
4660 : 00000;
4661 : 00000;
4662 : 00000;
4663 : 00000;
4664 : 00000;
4665 : 00000;
4666 : 00000;
4667 : 00000;
4670 : 00000;
4671 : 00000;
4672 : 00000;
4673 : 00000;
4674 : 00000;
4675 : 00000;
4676 : 00000;
4677 : 00000;
4700 : 00000;
4701 : 00000;
4702 : 00000;
4703 : 00000;
4704 : 00000;
4705 : 00000;
4706 : 00000;
4707 : 00000;
4710 : 00000;
4711 : 00000;
4712 : 00000;
4713 : 00000;
4714 : 00000;
4715 : 00000;
4716 : 00000;
4717 : 00000;
4720 : 00000;
4721 : 00000;
4722 : 00000;
4723 : 00000;
4724 : 00000;
4725 : 00000;
4726 : 00000;
4727 : 00000;
4730 : 00000;
4731 : 00000;
4732 : 00000;
4733 : 00000;
4734 : 00000;
4735 : 00000;
4736 : 00000;
4737 : 00000;
4740 : 00000;
4741 : 00000;
4742 : 00000;
4743 : 00000;
4744 : 00000;
4745 : 00000;
4746 : 00000;
4747 : 00000;
4750 : 00000;
4751 : 00000;
4752 : 00000;
4753 : 00000;
4754 : 00000;
4755 : 00000;
4756 : 00000;
4757 : 00000;
4760 : 00000;
4761 : 00000;
4762 : 00000;
4763 : 00000;
4764 : 00000;
4765 : 00000;
4766 : 00000;
4767 : 00000;
4770 : 00000;
4771 : 00000;
4772 : 00000;
4773 : 00000;
4774 : 00000;
4775 : 00000;
4776 : 00000;
4777 : 00000;
5000 : 00000;
5001 : 00000;
5002 : 00000;
5003 : 00000;
5004 : 00000;
5005 : 00000;
5006 : 00000;
5007 : 00000;
5010 : 00000;
5011 : 00000;
5012 : 00000;
5013 : 00000;
5014 : 00000;
5015 : 00000;
5016 : 00000;
5017 : 00000;
5020 : 00000;
5021 : 00000;
5022 : 00000;
5023 : 00000;
5024 : 00000;
5025 : 00000;
5026 : 00000;
5027 : 00000;
5030 : 00000;
5031 : 00000;
5032 : 00000;
5033 : 00000;
5034 : 00000;
5035 : 00000;
5036 : 00000;
5037 : 00000;
5040 : 00000;
5041 : 00000;
5042 : 00000;
5043 : 00000;
5044 : 00000;
5045 : 00000;
5046 : 00000;
5047 : 00000;
5050 : 00000;
5051 : 00000;
5052 : 00000;
5053 : 00000;
5054 : 00000;
5055 : 00000;
5056 : 00000;
5057 : 00000;
5060 : 00000;
5061 : 00000;
5062 : 00000;
5063 : 00000;
5064 : 00000;
5065 : 00000;
5066 : 00000;
5067 : 00000;
5070 : 00000;
5071 : 00000;
5072 : 00000;
5073 : 00000;
5074 : 00000;
5075 : 00000;
5076 : 00000;
5077 : 00000;
5100 : 00000;
5101 : 00000;
5102 : 00000;
5103 : 00000;
5104 : 00000;
5105 : 00000;
5106 : 00000;
5107 : 00000;
5110 : 00000;
5111 : 00000;
5112 : 00000;
5113 : 00000;
5114 : 00000;
5115 : 00000;
5116 : 00000;
5117 : 00000;
5120 : 00000;
5121 : 00000;
5122 : 00000;
5123 : 00000;
5124 : 00000;
5125 : 00000;
5126 : 00000;
5127 : 00000;
5130 : 00000;
5131 : 00000;
5132 : 00000;
5133 : 00000;
5134 : 00000;
5135 : 00000;
5136 : 00000;
5137 : 00000;
5140 : 00000;
5141 : 00000;
5142 : 00000;
5143 : 00000;
5144 : 00000;
5145 : 00000;
5146 : 00000;
5147 : 00000;
5150 : 00000;
5151 : 00000;
5152 : 00000;
5153 : 00000;
5154 : 00000;
5155 : 00000;
5156 : 00000;
5157 : 00000;
5160 : 00000;
5161 : 00000;
5162 : 00000;
5163 : 00000;
5164 : 00000;
5165 : 00000;
5166 : 00000;
5167 : 00000;
5170 : 00000;
5171 : 00000;
5172 : 00000;
5173 : 00000;
5174 : 00000;
5175 : 00000;
5176 : 00000;
5177 : 00000;
5200 : 00000;
5201 : 00000;
5202 : 00000;
5203 : 00000;
5204 : 00000;
5205 : 00000;
5206 : 00000;
5207 : 00000;
5210 : 00000;
5211 : 00000;
5212 : 00000;
5213 : 00000;
5214 : 00000;
5215 : 00000;
5216 : 00000;
5217 : 00000;
5220 : 00000;
5221 : 00000;
5222 : 00000;
5223 : 00000;
5224 : 00000;
5225 : 00000;
5226 : 00000;
5227 : 00000;
5230 : 00000;
5231 : 00000;
5232 : 00000;
5233 : 00000;
5234 : 00000;
5235 : 00000;
5236 : 00000;
5237 : 00000;
5240 : 00000;
5241 : 00000;
5242 : 00000;
5243 : 00000;
5244 : 00000;
5245 : 00000;
5246 : 00000;
5247 : 00000;
5250 : 00000;
5251 : 00000;
5252 : 00000;
5253 : 00000;
5254 : 00000;
5255 : 00000;
5256 : 00000;
5257 : 00000;
5260 : 00000;
5261 : 00000;
5262 : 00000;
5263 : 00000;
5264 : 00000;
5265 : 00000;
5266 : 00000;
5267 : 00000;
5270 : 00000;
5271 : 00000;
5272 : 00000;
5273 : 00000;
5274 : 00000;
5275 : 00000;
5276 : 00000;
5277 : 00000;
5300 : 00000;
5301 : 00000;
5302 : 00000;
5303 : 00000;
5304 : 00000;
5305 : 00000;
5306 : 00000;
5307 : 00000;
5310 : 00000;
5311 : 00000;
5312 : 00000;
5313 : 00000;
5314 : 00000;
5315 : 00000;
5316 : 00000;
5317 : 00000;
5320 : 00000;
5321 : 00000;
5322 : 00000;
5323 : 00000;
5324 : 00000;
5325 : 00000;
5326 : 00000;
5327 : 00000;
5330 : 00000;
5331 : 00000;
5332 : 00000;
5333 : 00000;
5334 : 00000;
5335 : 00000;
5336 : 00000;
5337 : 00000;
5340 : 00000;
5341 : 00000;
5342 : 00000;
5343 : 00000;
5344 : 00000;
5345 : 00000;
5346 : 00000;
5347 : 00000;
5350 : 00000;
5351 : 00000;
5352 : 00000;
5353 : 00000;
5354 : 00000;
5355 : 00000;
5356 : 00000;
5357 : 00000;
5360 : 00000;
5361 : 00000;
5362 : 00000;
5363 : 00000;
5364 : 00000;
5365 : 00000;
5366 : 00000;
5367 : 00000;
5370 : 00000;
5371 : 00000;
5372 : 00000;
5373 : 00000;
5374 : 00000;
5375 : 00000;
5376 : 00000;
5377 : 00000;
5400 : 00000;
5401 : 00000;
5402 : 00000;
5403 : 00000;
5404 : 00000;
5405 : 00000;
5406 : 00000;
5407 : 00000;
5410 : 00000;
5411 : 00000;
5412 : 00000;
5413 : 00000;
5414 : 00000;
5415 : 00000;
5416 : 00000;
5417 : 00000;
5420 : 00000;
5421 : 00000;
5422 : 00000;
5423 : 00000;
5424 : 00000;
5425 : 00000;
5426 : 00000;
5427 : 00000;
5430 : 00000;
5431 : 00000;
5432 : 00000;
5433 : 00000;
5434 : 00000;
5435 : 00000;
5436 : 00000;
5437 : 00000;
5440 : 00000;
5441 : 00000;
5442 : 00000;
5443 : 00000;
5444 : 00000;
5445 : 00000;
5446 : 00000;
5447 : 00000;
5450 : 00000;
5451 : 00000;
5452 : 00000;
5453 : 00000;
5454 : 00000;
5455 : 00000;
5456 : 00000;
5457 : 00000;
5460 : 00000;
5461 : 00000;
5462 : 00000;
5463 : 00000;
5464 : 00000;
5465 : 00000;
5466 : 00000;
5467 : 00000;
5470 : 00000;
5471 : 00000;
5472 : 00000;
5473 : 00000;
5474 : 00000;
5475 : 00000;
5476 : 00000;
5477 : 00000;
5500 : 00000;
5501 : 00000;
5502 : 00000;
5503 : 00000;
5504 : 00000;
5505 : 00000;
5506 : 00000;
5507 : 00000;
5510 : 00000;
5511 : 00000;
5512 : 00000;
5513 : 00000;
5514 : 00000;
5515 : 00000;
5516 : 00000;
5517 : 00000;
5520 : 00000;
5521 : 00000;
5522 : 00000;
5523 : 00000;
5524 : 00000;
5525 : 00000;
5526 : 00000;
5527 : 00000;
5530 : 00000;
5531 : 00000;
5532 : 00000;
5533 : 00000;
5534 : 00000;
5535 : 00000;
5536 : 00000;
5537 : 00000;
5540 : 00000;
5541 : 00000;
5542 : 00000;
5543 : 00000;
5544 : 00000;
5545 : 00000;
5546 : 00000;
5547 : 00000;
5550 : 00000;
5551 : 00000;
5552 : 00000;
5553 : 00000;
5554 : 00000;
5555 : 00000;
5556 : 00000;
5557 : 00000;
5560 : 00000;
5561 : 00000;
5562 : 00000;
5563 : 00000;
5564 : 00000;
5565 : 00000;
5566 : 00000;
5567 : 00000;
5570 : 00000;
5571 : 00000;
5572 : 00000;
5573 : 00000;
5574 : 00000;
5575 : 00000;
5576 : 00000;
5577 : 00000;
5600 : 00000;
5601 : 00000;
5602 : 00000;
5603 : 00000;
5604 : 00000;
5605 : 00000;
5606 : 00000;
5607 : 00000;
5610 : 00000;
5611 : 00000;
5612 : 00000;
5613 : 00000;
5614 : 00000;
5615 : 00000;
5616 : 00000;
5617 : 00000;
5620 : 00000;
5621 : 00000;
5622 : 00000;
5623 : 00000;
5624 : 00000;
5625 : 00000;
5626 : 00000;
5627 : 00000;
5630 : 00000;
5631 : 00000;
5632 : 00000;
5633 : 00000;
5634 : 00000;
5635 : 00000;
5636 : 00000;
5637 : 00000;
5640 : 00000;
5641 : 00000;
5642 : 00000;
5643 : 00000;
5644 : 00000;
5645 : 00000;
5646 : 00000;
5647 : 00000;
5650 : 00000;
5651 : 00000;
5652 : 00000;
5653 : 00000;
5654 : 00000;
5655 : 00000;
5656 : 00000;
5657 : 00000;
5660 : 00000;
5661 : 00000;
5662 : 00000;
5663 : 00000;
5664 : 00000;
5665 : 00000;
5666 : 00000;
5667 : 00000;
5670 : 00000;
5671 : 00000;
5672 : 00000;
5673 : 00000;
5674 : 00000;
5675 : 00000;
5676 : 00000;
5677 : 00000;
5700 : 00000;
5701 : 00000;
5702 : 00000;
5703 : 00000;
5704 : 00000;
5705 : 00000;
5706 : 00000;
5707 : 00000;
5710 : 00000;
5711 : 00000;
5712 : 00000;
5713 : 00000;
5714 : 00000;
5715 : 00000;
5716 : 00000;
5717 : 00000;
5720 : 00000;
5721 : 00000;
5722 : 00000;
5723 : 00000;
5724 : 00000;
5725 : 00000;
5726 : 00000;
5727 : 00000;
5730 : 00000;
5731 : 00000;
5732 : 00000;
5733 : 00000;
5734 : 00000;
5735 : 00000;
5736 : 00000;
5737 : 00000;
5740 : 00000;
5741 : 00000;
5742 : 00000;
5743 : 00000;
5744 : 00000;
5745 : 00000;
5746 : 00000;
5747 : 00000;
5750 : 00000;
5751 : 00000;
5752 : 00000;
5753 : 00000;
5754 : 00000;
5755 : 00000;
5756 : 00000;
5757 : 00000;
5760 : 00000;
5761 : 00000;
5762 : 00000;
5763 : 00000;
5764 : 00000;
5765 : 00000;
5766 : 00000;
5767 : 00000;
5770 : 00000;
5771 : 00000;
5772 : 00000;
5773 : 00000;
5774 : 00000;
5775 : 00000;
5776 : 00000;
5777 : 00000;
6000 : 00000;
6001 : 00000;
6002 : 00000;
6003 : 00000;
6004 : 00000;
6005 : 00000;
6006 : 00000;
6007 : 00000;
6010 : 00000;
6011 : 00000;
6012 : 00000;
6013 : 00000;
6014 : 00000;
6015 : 00000;
6016 : 00000;
6017 : 00000;
6020 : 00000;
6021 : 00000;
6022 : 00000;
6023 : 00000;
6024 : 00000;
6025 : 00000;
6026 : 00000;
6027 : 00000;
6030 : 00000;
6031 : 00000;
6032 : 00000;
6033 : 00000;
6034 : 00000;
6035 : 00000;
6036 : 00000;
6037 : 00000;
6040 : 00000;
6041 : 00000;
6042 : 00000;
6043 : 00000;
6044 : 00000;
6045 : 00000;
6046 : 00000;
6047 : 00000;
6050 : 00000;
6051 : 00000;
6052 : 00000;
6053 : 00000;
6054 : 00000;
6055 : 00000;
6056 : 00000;
6057 : 00000;
6060 : 00000;
6061 : 00000;
6062 : 00000;
6063 : 00000;
6064 : 00000;
6065 : 00000;
6066 : 00000;
6067 : 00000;
6070 : 00000;
6071 : 00000;
6072 : 00000;
6073 : 00000;
6074 : 00000;
6075 : 00000;
6076 : 00000;
6077 : 00000;
6100 : 00000;
6101 : 00000;
6102 : 00000;
6103 : 00000;
6104 : 00000;
6105 : 00000;
6106 : 00000;
6107 : 00000;
6110 : 00000;
6111 : 00000;
6112 : 00000;
6113 : 00000;
6114 : 00000;
6115 : 00000;
6116 : 00000;
6117 : 00000;
6120 : 00000;
6121 : 00000;
6122 : 00000;
6123 : 00000;
6124 : 00000;
6125 : 00000;
6126 : 00000;
6127 : 00000;
6130 : 00000;
6131 : 00000;
6132 : 00000;
6133 : 00000;
6134 : 00000;
6135 : 00000;
6136 : 00000;
6137 : 00000;
6140 : 00000;
6141 : 00000;
6142 : 00000;
6143 : 00000;
6144 : 00000;
6145 : 00000;
6146 : 00000;
6147 : 00000;
6150 : 00000;
6151 : 00000;
6152 : 00000;
6153 : 00000;
6154 : 00000;
6155 : 00000;
6156 : 00000;
6157 : 00000;
6160 : 00000;
6161 : 00000;
6162 : 00000;
6163 : 00000;
6164 : 00000;
6165 : 00000;
6166 : 00000;
6167 : 00000;
6170 : 00000;
6171 : 00000;
6172 : 00000;
6173 : 00000;
6174 : 00000;
6175 : 00000;
6176 : 00000;
6177 : 00000;
6200 : 00000;
6201 : 00000;
6202 : 00000;
6203 : 00000;
6204 : 00000;
6205 : 00000;
6206 : 00000;
6207 : 00000;
6210 : 00000;
6211 : 00000;
6212 : 00000;
6213 : 00000;
6214 : 00000;
6215 : 00000;
6216 : 00000;
6217 : 00000;
6220 : 00000;
6221 : 00000;
6222 : 00000;
6223 : 00000;
6224 : 00000;
6225 : 00000;
6226 : 00000;
6227 : 00000;
6230 : 00000;
6231 : 00000;
6232 : 00000;
6233 : 00000;
6234 : 00000;
6235 : 00000;
6236 : 00000;
6237 : 00000;
6240 : 00000;
6241 : 00000;
6242 : 00000;
6243 : 00000;
6244 : 00000;
6245 : 00000;
6246 : 00000;
6247 : 00000;
6250 : 00000;
6251 : 00000;
6252 : 00000;
6253 : 00000;
6254 : 00000;
6255 : 00000;
6256 : 00000;
6257 : 00000;
6260 : 00000;
6261 : 00000;
6262 : 00000;
6263 : 00000;
6264 : 00000;
6265 : 00000;
6266 : 00000;
6267 : 00000;
6270 : 00000;
6271 : 00000;
6272 : 00000;
6273 : 00000;
6274 : 00000;
6275 : 00000;
6276 : 00000;
6277 : 00000;
6300 : 00000;
6301 : 00000;
6302 : 00000;
6303 : 00000;
6304 : 00000;
6305 : 00000;
6306 : 00000;
6307 : 00000;
6310 : 00000;
6311 : 00000;
6312 : 00000;
6313 : 00000;
6314 : 00000;
6315 : 00000;
6316 : 00000;
6317 : 00000;
6320 : 00000;
6321 : 00000;
6322 : 00000;
6323 : 00000;
6324 : 00000;
6325 : 00000;
6326 : 00000;
6327 : 00000;
6330 : 00000;
6331 : 00000;
6332 : 00000;
6333 : 00000;
6334 : 00000;
6335 : 00000;
6336 : 00000;
6337 : 00000;
6340 : 00000;
6341 : 00000;
6342 : 00000;
6343 : 00000;
6344 : 00000;
6345 : 00000;
6346 : 00000;
6347 : 00000;
6350 : 00000;
6351 : 00000;
6352 : 00000;
6353 : 00000;
6354 : 00000;
6355 : 00000;
6356 : 00000;
6357 : 00000;
6360 : 00000;
6361 : 00000;
6362 : 00000;
6363 : 00000;
6364 : 00000;
6365 : 00000;
6366 : 00000;
6367 : 00000;
6370 : 00000;
6371 : 00000;
6372 : 00000;
6373 : 00000;
6374 : 00000;
6375 : 00000;
6376 : 00000;
6377 : 00000;
6400 : 00000;
6401 : 00000;
6402 : 00000;
6403 : 00000;
6404 : 00000;
6405 : 00000;
6406 : 00000;
6407 : 00000;
6410 : 00000;
6411 : 00000;
6412 : 00000;
6413 : 00000;
6414 : 00000;
6415 : 00000;
6416 : 00000;
6417 : 00000;
6420 : 00000;
6421 : 00000;
6422 : 00000;
6423 : 00000;
6424 : 00000;
6425 : 00000;
6426 : 00000;
6427 : 00000;
6430 : 00000;
6431 : 00000;
6432 : 00000;
6433 : 00000;
6434 : 00000;
6435 : 00000;
6436 : 00000;
6437 : 00000;
6440 : 00000;
6441 : 00000;
6442 : 00000;
6443 : 00000;
6444 : 00000;
6445 : 00000;
6446 : 00000;
6447 : 00000;
6450 : 00000;
6451 : 00000;
6452 : 00000;
6453 : 00000;
6454 : 00000;
6455 : 00000;
6456 : 00000;
6457 : 00000;
6460 : 00000;
6461 : 00000;
6462 : 00000;
6463 : 00000;
6464 : 00000;
6465 : 00000;
6466 : 00000;
6467 : 00000;
6470 : 00000;
6471 : 00000;
6472 : 00000;
6473 : 00000;
6474 : 00000;
6475 : 00000;
6476 : 00000;
6477 : 00000;
6500 : 00000;
6501 : 00000;
6502 : 00000;
6503 : 00000;
6504 : 00000;
6505 : 00000;
6506 : 00000;
6507 : 00000;
6510 : 00000;
6511 : 00000;
6512 : 00000;
6513 : 00000;
6514 : 00000;
6515 : 00000;
6516 : 00000;
6517 : 00000;
6520 : 00000;
6521 : 00000;
6522 : 00000;
6523 : 00000;
6524 : 00000;
6525 : 00000;
6526 : 00000;
6527 : 00000;
6530 : 00000;
6531 : 00000;
6532 : 00000;
6533 : 00000;
6534 : 00000;
6535 : 00000;
6536 : 00000;
6537 : 00000;
6540 : 00000;
6541 : 00000;
6542 : 00000;
6543 : 00000;
6544 : 00000;
6545 : 00000;
6546 : 00000;
6547 : 00000;
6550 : 00000;
6551 : 00000;
6552 : 00000;
6553 : 00000;
6554 : 00000;
6555 : 00000;
6556 : 00000;
6557 : 00000;
6560 : 00000;
6561 : 00000;
6562 : 00000;
6563 : 00000;
6564 : 00000;
6565 : 00000;
6566 : 00000;
6567 : 00000;
6570 : 00000;
6571 : 00000;
6572 : 00000;
6573 : 00000;
6574 : 00000;
6575 : 00000;
6576 : 00000;
6577 : 00000;
6600 : 00000;
6601 : 00000;
6602 : 00000;
6603 : 00000;
6604 : 00000;
6605 : 00000;
6606 : 00000;
6607 : 00000;
6610 : 00000;
6611 : 00000;
6612 : 00000;
6613 : 00000;
6614 : 00000;
6615 : 00000;
6616 : 00000;
6617 : 00000;
6620 : 00000;
6621 : 00000;
6622 : 00000;
6623 : 00000;
6624 : 00000;
6625 : 00000;
6626 : 00000;
6627 : 00000;
6630 : 00000;
6631 : 00000;
6632 : 00000;
6633 : 00000;
6634 : 00000;
6635 : 00000;
6636 : 00000;
6637 : 00000;
6640 : 00000;
6641 : 00000;
6642 : 00000;
6643 : 00000;
6644 : 00000;
6645 : 00000;
6646 : 00000;
6647 : 00000;
6650 : 00000;
6651 : 00000;
6652 : 00000;
6653 : 00000;
6654 : 00000;
6655 : 00000;
6656 : 00000;
6657 : 00000;
6660 : 00000;
6661 : 00000;
6662 : 00000;
6663 : 00000;
6664 : 00000;
6665 : 00000;
6666 : 00000;
6667 : 00000;
6670 : 00000;
6671 : 00000;
6672 : 00000;
6673 : 00000;
6674 : 00000;
6675 : 00000;
6676 : 00000;
6677 : 00000;
6700 : 00000;
6701 : 00000;
6702 : 00000;
6703 : 00000;
6704 : 00000;
6705 : 00000;
6706 : 00000;
6707 : 00000;
6710 : 00000;
6711 : 00000;
6712 : 00000;
6713 : 00000;
6714 : 00000;
6715 : 00000;
6716 : 00000;
6717 : 00000;
6720 : 00000;
6721 : 00000;
6722 : 00000;
6723 : 00000;
6724 : 00000;
6725 : 00000;
6726 : 00000;
6727 : 00000;
6730 : 00000;
6731 : 00000;
6732 : 00000;
6733 : 00000;
6734 : 00000;
6735 : 00000;
6736 : 00000;
6737 : 00000;
6740 : 00000;
6741 : 00000;
6742 : 00000;
6743 : 00000;
6744 : 00000;
6745 : 00000;
6746 : 00000;
6747 : 00000;
6750 : 00000;
6751 : 00000;
6752 : 00000;
6753 : 00000;
6754 : 00000;
6755 : 00000;
6756 : 00000;
6757 : 00000;
6760 : 00000;
6761 : 00000;
6762 : 00000;
6763 : 00000;
6764 : 00000;
6765 : 00000;
6766 : 00000;
6767 : 00000;
6770 : 00000;
6771 : 00000;
6772 : 00000;
6773 : 00000;
6774 : 00000;
6775 : 00000;
6776 : 00000;
6777 : 00000;
7000 : 00000;
7001 : 00000;
7002 : 00000;
7003 : 00000;
7004 : 00000;
7005 : 00000;
7006 : 00000;
7007 : 00000;
7010 : 00000;
7011 : 00000;
7012 : 00000;
7013 : 00000;
7014 : 00000;
7015 : 00000;
7016 : 00000;
7017 : 00000;
7020 : 00000;
7021 : 00000;
7022 : 00000;
7023 : 00000;
7024 : 00000;
7025 : 00000;
7026 : 00000;
7027 : 00000;
7030 : 00000;
7031 : 00000;
7032 : 00000;
7033 : 00000;
7034 : 00000;
7035 : 00000;
7036 : 00000;
7037 : 00000;
7040 : 00000;
7041 : 00000;
7042 : 00000;
7043 : 00000;
7044 : 00000;
7045 : 00000;
7046 : 00000;
7047 : 00000;
7050 : 00000;
7051 : 00000;
7052 : 00000;
7053 : 00000;
7054 : 00000;
7055 : 00000;
7056 : 00000;
7057 : 00000;
7060 : 00000;
7061 : 00000;
7062 : 00000;
7063 : 00000;
7064 : 00000;
7065 : 00000;
7066 : 00000;
7067 : 00000;
7070 : 00000;
7071 : 00000;
7072 : 00000;
7073 : 00000;
7074 : 00000;
7075 : 00000;
7076 : 00000;
7077 : 00000;
7100 : 00000;
7101 : 00000;
7102 : 00000;
7103 : 00000;
7104 : 00000;
7105 : 00000;
7106 : 00000;
7107 : 00000;
7110 : 00000;
7111 : 00000;
7112 : 00000;
7113 : 00000;
7114 : 00000;
7115 : 00000;
7116 : 00000;
7117 : 00000;
7120 : 00000;
7121 : 00000;
7122 : 00000;
7123 : 00000;
7124 : 00000;
7125 : 00000;
7126 : 00000;
7127 : 00000;
7130 : 00000;
7131 : 00000;
7132 : 00000;
7133 : 00000;
7134 : 00000;
7135 : 00000;
7136 : 00000;
7137 : 00000;
7140 : 00000;
7141 : 00000;
7142 : 00000;
7143 : 00000;
7144 : 00000;
7145 : 00000;
7146 : 00000;
7147 : 00000;
7150 : 00000;
7151 : 00000;
7152 : 00000;
7153 : 00000;
7154 : 00000;
7155 : 00000;
7156 : 00000;
7157 : 00000;
7160 : 00000;
7161 : 00000;
7162 : 00000;
7163 : 00000;
7164 : 00000;
7165 : 00000;
7166 : 00000;
7167 : 00000;
7170 : 00000;
7171 : 00000;
7172 : 00000;
7173 : 00000;
7174 : 00000;
7175 : 00000;
7176 : 00000;
7177 : 00000;
7200 : 00000;
7201 : 00000;
7202 : 00000;
7203 : 00000;
7204 : 00000;
7205 : 00000;
7206 : 00000;
7207 : 00000;
7210 : 00000;
7211 : 00000;
7212 : 00000;
7213 : 00000;
7214 : 00000;
7215 : 00000;
7216 : 00000;
7217 : 00000;
7220 : 00000;
7221 : 00000;
7222 : 00000;
7223 : 00000;
7224 : 00000;
7225 : 00000;
7226 : 00000;
7227 : 00000;
7230 : 00000;
7231 : 00000;
7232 : 00000;
7233 : 00000;
7234 : 00000;
7235 : 00000;
7236 : 00000;
7237 : 00000;
7240 : 00000;
7241 : 00000;
7242 : 00000;
7243 : 00000;
7244 : 00000;
7245 : 00000;
7246 : 00000;
7247 : 00000;
7250 : 00000;
7251 : 00000;
7252 : 00000;
7253 : 00000;
7254 : 00000;
7255 : 00000;
7256 : 00000;
7257 : 00000;
7260 : 00000;
7261 : 00000;
7262 : 00000;
7263 : 00000;
7264 : 00000;
7265 : 00000;
7266 : 00000;
7267 : 00000;
7270 : 00000;
7271 : 00000;
7272 : 00000;
7273 : 00000;
7274 : 00000;
7275 : 00000;
7276 : 00000;
7277 : 00000;
7300 : 00000;
7301 : 00000;
7302 : 00000;
7303 : 00000;
7304 : 00000;
7305 : 00000;
7306 : 00000;
7307 : 00000;
7310 : 00000;
7311 : 00000;
7312 : 00000;
7313 : 00000;
7314 : 00000;
7315 : 00000;
7316 : 00000;
7317 : 00000;
7320 : 00000;
7321 : 00000;
7322 : 00000;
7323 : 00000;
7324 : 00000;
7325 : 00000;
7326 : 00000;
7327 : 00000;
7330 : 00000;
7331 : 00000;
7332 : 00000;
7333 : 00000;
7334 : 00000;
7335 : 00000;
7336 : 00000;
7337 : 00000;
7340 : 00000;
7341 : 00000;
7342 : 00000;
7343 : 00000;
7344 : 00000;
7345 : 00000;
7346 : 00000;
7347 : 00000;
7350 : 00000;
7351 : 00000;
7352 : 00000;
7353 : 00000;
7354 : 00000;
7355 : 00000;
7356 : 00000;
7357 : 00000;
7360 : 00000;
7361 : 00000;
7362 : 00000;
7363 : 00000;
7364 : 00000;
7365 : 00000;
7366 : 00000;
7367 : 00000;
7370 : 00000;
7371 : 00000;
7372 : 00000;
7373 : 00000;
7374 : 00000;
7375 : 00000;
7376 : 00000;
7377 : 00000;
7400 : 00000;
7401 : 00000;
7402 : 00000;
7403 : 00000;
7404 : 00000;
7405 : 00000;
7406 : 00000;
7407 : 00000;
7410 : 00000;
7411 : 00000;
7412 : 00000;
7413 : 00000;
7414 : 00000;
7415 : 00000;
7416 : 00000;
7417 : 00000;
7420 : 00000;
7421 : 00000;
7422 : 00000;
7423 : 00000;
7424 : 00000;
7425 : 00000;
7426 : 00000;
7427 : 00000;
7430 : 00000;
7431 : 00000;
7432 : 00000;
7433 : 00000;
7434 : 00000;
7435 : 00000;
7436 : 00000;
7437 : 00000;
7440 : 00000;
7441 : 00000;
7442 : 00000;
7443 : 00000;
7444 : 00000;
7445 : 00000;
7446 : 00000;
7447 : 00000;
7450 : 00000;
7451 : 00000;
7452 : 00000;
7453 : 00000;
7454 : 00000;
7455 : 00000;
7456 : 00000;
7457 : 00000;
7460 : 00000;
7461 : 00000;
7462 : 00000;
7463 : 00000;
7464 : 00000;
7465 : 00000;
7466 : 00000;
7467 : 00000;
7470 : 00000;
7471 : 00000;
7472 : 00000;
7473 : 00000;
7474 : 00000;
7475 : 00000;
7476 : 00000;
7477 : 00000;
7500 : 00000;
7501 : 00000;
7502 : 00000;
7503 : 00000;
7504 : 00000;
7505 : 00000;
7506 : 00000;
7507 : 00000;
7510 : 00000;
7511 : 00000;
7512 : 00000;
7513 : 00000;
7514 : 00000;
7515 : 00000;
7516 : 00000;
7517 : 00000;
7520 : 00000;
7521 : 00000;
7522 : 00000;
7523 : 00000;
7524 : 00000;
7525 : 00000;
7526 : 00000;
7527 : 00000;
7530 : 00000;
7531 : 00000;
7532 : 00000;
7533 : 00000;
7534 : 00000;
7535 : 00000;
7536 : 00000;
7537 : 00000;
7540 : 00000;
7541 : 00000;
7542 : 00000;
7543 : 00000;
7544 : 00000;
7545 : 00000;
7546 : 00000;
7547 : 00000;
7550 : 00000;
7551 : 00000;
7552 : 00000;
7553 : 00000;
7554 : 00000;
7555 : 00000;
7556 : 00000;
7557 : 00000;
7560 : 00000;
7561 : 00000;
7562 : 00000;
7563 : 00000;
7564 : 00000;
7565 : 00000;
7566 : 00000;
7567 : 00000;
7570 : 00000;
7571 : 00000;
7572 : 00000;
7573 : 00000;
7574 : 00000;
7575 : 00000;
7576 : 00000;
7577 : 00000;
7600 : 00000;
7601 : 00000;
7602 : 00000;
7603 : 00000;
7604 : 00000;
7605 : 00000;
7606 : 00000;
7607 : 00000;
7610 : 00000;
7611 : 00000;
7612 : 00000;
7613 : 00000;
7614 : 00000;
7615 : 00000;
7616 : 00000;
7617 : 00000;
7620 : 00000;
7621 : 00000;
7622 : 00000;
7623 : 00000;
7624 : 00000;
7625 : 00000;
7626 : 00000;
7627 : 00000;
7630 : 00000;
7631 : 00000;
7632 : 00000;
7633 : 00000;
7634 : 00000;
7635 : 00000;
7636 : 00000;
7637 : 00000;
7640 : 00000;
7641 : 00000;
7642 : 00000;
7643 : 00000;
7644 : 00000;
7645 : 00000;
7646 : 00000;
7647 : 00000;
7650 : 00000;
7651 : 00000;
7652 : 00000;
7653 : 00000;
7654 : 00000;
7655 : 00000;
7656 : 00000;
7657 : 00000;
7660 : 00000;
7661 : 00000;
7662 : 00000;
7663 : 00000;
7664 : 00000;
7665 : 00000;
7666 : 00000;
7667 : 00000;
7670 : 00000;
7671 : 00000;
7672 : 00000;
7673 : 00000;
7674 : 00000;
7675 : 00000;
7676 : 00000;
7677 : 00000;
7700 : 00000;
7701 : 00000;
7702 : 00000;
7703 : 00000;
7704 : 00000;
7705 : 00000;
7706 : 00000;
7707 : 00000;
7710 : 00000;
7711 : 00000;
7712 : 00000;
7713 : 00000;
7714 : 00000;
7715 : 00000;
7716 : 00000;
7717 : 00000;
7720 : 00000;
7721 : 00000;
7722 : 00000;
7723 : 00000;
7724 : 00000;
7725 : 00000;
7726 : 00000;
7727 : 00000;
7730 : 00000;
7731 : 00000;
7732 : 00000;
7733 : 00000;
7734 : 00000;
7735 : 00000;
7736 : 00000;
7737 : 00000;
7740 : 00000;
7741 : 00000;
7742 : 00000;
7743 : 00000;
7744 : 00000;
7745 : 00000;
7746 : 00000;
7747 : 00000;
7750 : 00000;
7751 : 00000;
7752 : 00000;
7753 : 00000;
7754 : 00000;
7755 : 00000;
7756 : 00000;
7757 : 00000;
7760 : 00000;
7761 : 00000;
7762 : 00000;
7763 : 00000;
7764 : 00000;
7765 : 00000;
7766 : 00000;
7767 : 00000;
7770 : 00000;
7771 : 00000;
7772 : 00000;
7773 : 00000;
7774 : 00000;
7775 : 00000;
7776 : 00000;
7777 : 00000;
10000 : 00000;
10001 : 00000;
10002 : 00000;
10003 : 00000;
10004 : 00000;
10005 : 00000;
10006 : 00000;
10007 : 00000;
10010 : 00000;
10011 : 00000;
10012 : 00000;
10013 : 00000;
10014 : 00000;
10015 : 00000;
10016 : 00000;
10017 : 00000;
10020 : 00000;
10021 : 00000;
10022 : 00000;
10023 : 00000;
10024 : 00000;
10025 : 00000;
10026 : 00000;
10027 : 00000;
10030 : 00000;
10031 : 00000;
10032 : 00000;
10033 : 00000;
10034 : 00000;
10035 : 00000;
10036 : 00000;
10037 : 00000;
10040 : 00000;
10041 : 00000;
10042 : 00000;
10043 : 00000;
10044 : 00000;
10045 : 00000;
10046 : 00000;
10047 : 00000;
10050 : 00000;
10051 : 00000;
10052 : 00000;
10053 : 00000;
10054 : 00000;
10055 : 00000;
10056 : 00000;
10057 : 00000;
10060 : 00000;
10061 : 00000;
10062 : 00000;
10063 : 00000;
10064 : 00000;
10065 : 00000;
10066 : 00000;
10067 : 00000;
10070 : 00000;
10071 : 00000;
10072 : 00000;
10073 : 00000;
10074 : 04074;
10075 : 04075;
10076 : 67610;
10077 : 00000;
10100 : 00000;
10101 : 00000;
10102 : 00000;
10103 : 00000;
10104 : 00000;
10105 : 00000;
10106 : 00000;
10107 : 00000;
10110 : 00000;
10111 : 00000;
10112 : 00000;
10113 : 00000;
10114 : 00000;
10115 : 00000;
10116 : 00000;
10117 : 00000;
10120 : 00000;
10121 : 00000;
10122 : 00000;
10123 : 00000;
10124 : 00000;
10125 : 00000;
10126 : 00000;
10127 : 00000;
10130 : 00000;
10131 : 00000;
10132 : 00000;
10133 : 00000;
10134 : 00000;
10135 : 00000;
10136 : 00000;
10137 : 00000;
10140 : 00000;
10141 : 00000;
10142 : 00000;
10143 : 00000;
10144 : 00000;
10145 : 00000;
10146 : 00000;
10147 : 00000;
10150 : 00000;
10151 : 00000;
10152 : 00000;
10153 : 00000;
10154 : 00000;
10155 : 00000;
10156 : 00000;
10157 : 00000;
10160 : 00000;
10161 : 00000;
10162 : 00000;
10163 : 00000;
10164 : 00000;
10165 : 00000;
10166 : 00000;
10167 : 00000;
10170 : 00000;
10171 : 00000;
10172 : 00000;
10173 : 00000;
10174 : 00000;
10175 : 00000;
10176 : 00000;
10177 : 00000;
10200 : 00000;
10201 : 00000;
10202 : 00000;
10203 : 00000;
10204 : 00000;
10205 : 00000;
10206 : 00000;
10207 : 00000;
10210 : 00000;
10211 : 00000;
10212 : 00000;
10213 : 00000;
10214 : 00000;
10215 : 00000;
10216 : 00000;
10217 : 00000;
10220 : 00000;
10221 : 00000;
10222 : 00000;
10223 : 00000;
10224 : 00000;
10225 : 00000;
10226 : 00000;
10227 : 00000;
10230 : 00000;
10231 : 00000;
10232 : 00000;
10233 : 00000;
10234 : 00000;
10235 : 00000;
10236 : 00000;
10237 : 00000;
10240 : 00000;
10241 : 00000;
10242 : 00000;
10243 : 00000;
10244 : 00000;
10245 : 00000;
10246 : 00000;
10247 : 00000;
10250 : 00000;
10251 : 00000;
10252 : 00000;
10253 : 00000;
10254 : 00000;
10255 : 00000;
10256 : 00000;
10257 : 00000;
10260 : 00000;
10261 : 00000;
10262 : 00000;
10263 : 00000;
10264 : 00000;
10265 : 00000;
10266 : 00000;
10267 : 00000;
10270 : 00000;
10271 : 00000;
10272 : 00000;
10273 : 00000;
10274 : 00000;
10275 : 00000;
10276 : 00000;
10277 : 00000;
10300 : 00000;
10301 : 00000;
10302 : 00000;
10303 : 00000;
10304 : 00000;
10305 : 00000;
10306 : 00000;
10307 : 00000;
10310 : 00000;
10311 : 00000;
10312 : 00000;
10313 : 00000;
10314 : 00000;
10315 : 00000;
10316 : 00000;
10317 : 00000;
10320 : 00000;
10321 : 00000;
10322 : 00000;
10323 : 00000;
10324 : 00000;
10325 : 00000;
10326 : 00000;
10327 : 00000;
10330 : 00000;
10331 : 00000;
10332 : 00000;
10333 : 00000;
10334 : 00000;
10335 : 00000;
10336 : 00000;
10337 : 00000;
10340 : 00000;
10341 : 00000;
10342 : 00000;
10343 : 00000;
10344 : 00000;
10345 : 00000;
10346 : 00000;
10347 : 00000;
10350 : 00000;
10351 : 00000;
10352 : 00000;
10353 : 00000;
10354 : 00000;
10355 : 00000;
10356 : 00000;
10357 : 00000;
10360 : 00000;
10361 : 00000;
10362 : 00000;
10363 : 00000;
10364 : 00000;
10365 : 00000;
10366 : 00000;
10367 : 00000;
10370 : 00000;
10371 : 00000;
10372 : 00000;
10373 : 00000;
10374 : 00000;
10375 : 00000;
10376 : 00000;
10377 : 00000;
10400 : 00000;
10401 : 00000;
10402 : 00000;
10403 : 00000;
10404 : 00000;
10405 : 00000;
10406 : 00000;
10407 : 00000;
10410 : 00000;
10411 : 00000;
10412 : 00000;
10413 : 00000;
10414 : 00000;
10415 : 00000;
10416 : 00000;
10417 : 00000;
10420 : 00000;
10421 : 00000;
10422 : 00000;
10423 : 00000;
10424 : 00000;
10425 : 00000;
10426 : 00000;
10427 : 00000;
10430 : 00000;
10431 : 00000;
10432 : 00000;
10433 : 00000;
10434 : 00000;
10435 : 00000;
10436 : 00000;
10437 : 00000;
10440 : 00000;
10441 : 00000;
10442 : 00000;
10443 : 00000;
10444 : 00000;
10445 : 00000;
10446 : 00000;
10447 : 00000;
10450 : 00000;
10451 : 00000;
10452 : 00000;
10453 : 00000;
10454 : 00000;
10455 : 00000;
10456 : 00000;
10457 : 00000;
10460 : 00000;
10461 : 00000;
10462 : 00000;
10463 : 00000;
10464 : 00000;
10465 : 00000;
10466 : 00000;
10467 : 00000;
10470 : 00000;
10471 : 00000;
10472 : 00000;
10473 : 00000;
10474 : 00000;
10475 : 00000;
10476 : 00000;
10477 : 00000;
10500 : 00000;
10501 : 00000;
10502 : 00000;
10503 : 00000;
10504 : 00000;
10505 : 00000;
10506 : 00000;
10507 : 00000;
10510 : 00000;
10511 : 00000;
10512 : 00000;
10513 : 00000;
10514 : 00000;
10515 : 00000;
10516 : 00000;
10517 : 00000;
10520 : 00000;
10521 : 00000;
10522 : 00000;
10523 : 00000;
10524 : 00000;
10525 : 00000;
10526 : 00000;
10527 : 00000;
10530 : 00000;
10531 : 00000;
10532 : 00000;
10533 : 00000;
10534 : 00000;
10535 : 00000;
10536 : 00000;
10537 : 00000;
10540 : 00000;
10541 : 00000;
10542 : 00000;
10543 : 00000;
10544 : 00000;
10545 : 00000;
10546 : 00000;
10547 : 00000;
10550 : 00000;
10551 : 00000;
10552 : 00000;
10553 : 00000;
10554 : 00000;
10555 : 00000;
10556 : 00000;
10557 : 00000;
10560 : 00000;
10561 : 00000;
10562 : 00000;
10563 : 00000;
10564 : 00000;
10565 : 00000;
10566 : 00000;
10567 : 00000;
10570 : 00000;
10571 : 00000;
10572 : 00000;
10573 : 00000;
10574 : 00000;
10575 : 00000;
10576 : 00000;
10577 : 00000;
10600 : 00000;
10601 : 00000;
10602 : 00000;
10603 : 00000;
10604 : 00000;
10605 : 00000;
10606 : 00000;
10607 : 00000;
10610 : 00000;
10611 : 00000;
10612 : 00000;
10613 : 00000;
10614 : 00000;
10615 : 00000;
10616 : 00000;
10617 : 00000;
10620 : 00000;
10621 : 00000;
10622 : 00000;
10623 : 00000;
10624 : 00000;
10625 : 00000;
10626 : 00000;
10627 : 00000;
10630 : 00000;
10631 : 00000;
10632 : 00000;
10633 : 00000;
10634 : 00000;
10635 : 00000;
10636 : 00000;
10637 : 00000;
10640 : 00000;
10641 : 00000;
10642 : 00000;
10643 : 00000;
10644 : 00000;
10645 : 00000;
10646 : 00000;
10647 : 00000;
10650 : 00000;
10651 : 00000;
10652 : 00000;
10653 : 00000;
10654 : 00000;
10655 : 00000;
10656 : 00000;
10657 : 00000;
10660 : 00000;
10661 : 00000;
10662 : 00000;
10663 : 00000;
10664 : 00000;
10665 : 00000;
10666 : 00000;
10667 : 00000;
10670 : 00000;
10671 : 00000;
10672 : 00000;
10673 : 00000;
10674 : 00000;
10675 : 00000;
10676 : 00000;
10677 : 00000;
10700 : 00000;
10701 : 00000;
10702 : 00000;
10703 : 00000;
10704 : 00000;
10705 : 00000;
10706 : 00000;
10707 : 00000;
10710 : 00000;
10711 : 00000;
10712 : 00000;
10713 : 00000;
10714 : 00000;
10715 : 00000;
10716 : 00000;
10717 : 00000;
10720 : 00000;
10721 : 00000;
10722 : 00000;
10723 : 00000;
10724 : 00000;
10725 : 00000;
10726 : 00000;
10727 : 00000;
10730 : 00000;
10731 : 00000;
10732 : 00000;
10733 : 00000;
10734 : 00000;
10735 : 00000;
10736 : 00000;
10737 : 00000;
10740 : 00000;
10741 : 00000;
10742 : 00000;
10743 : 00000;
10744 : 00000;
10745 : 00000;
10746 : 00000;
10747 : 00000;
10750 : 00000;
10751 : 00000;
10752 : 00000;
10753 : 00000;
10754 : 00000;
10755 : 00000;
10756 : 00000;
10757 : 00000;
10760 : 00000;
10761 : 00000;
10762 : 00000;
10763 : 00000;
10764 : 00000;
10765 : 00000;
10766 : 00000;
10767 : 00000;
10770 : 00000;
10771 : 00000;
10772 : 00000;
10773 : 00000;
10774 : 00000;
10775 : 00000;
10776 : 00000;
10777 : 00000;
11000 : 00000;
11001 : 00000;
11002 : 00000;
11003 : 00000;
11004 : 00000;
11005 : 00000;
11006 : 00000;
11007 : 00000;
11010 : 00000;
11011 : 00000;
11012 : 00000;
11013 : 00000;
11014 : 00000;
11015 : 00000;
11016 : 00000;
11017 : 00000;
11020 : 00000;
11021 : 00000;
11022 : 00000;
11023 : 00000;
11024 : 00000;
11025 : 00000;
11026 : 00000;
11027 : 00000;
11030 : 00000;
11031 : 00000;
11032 : 00000;
11033 : 00000;
11034 : 00000;
11035 : 00000;
11036 : 00000;
11037 : 00000;
11040 : 00000;
11041 : 00000;
11042 : 00000;
11043 : 00000;
11044 : 00000;
11045 : 00000;
11046 : 00000;
11047 : 00000;
11050 : 00000;
11051 : 00000;
11052 : 00000;
11053 : 00000;
11054 : 00000;
11055 : 00000;
11056 : 00000;
11057 : 00000;
11060 : 00000;
11061 : 00000;
11062 : 00000;
11063 : 00000;
11064 : 00000;
11065 : 00000;
11066 : 00000;
11067 : 00000;
11070 : 00000;
11071 : 00000;
11072 : 00000;
11073 : 00000;
11074 : 00000;
11075 : 00000;
11076 : 00000;
11077 : 00000;
11100 : 00000;
11101 : 00000;
11102 : 00000;
11103 : 00000;
11104 : 00000;
11105 : 00000;
11106 : 00000;
11107 : 00000;
11110 : 00000;
11111 : 00000;
11112 : 00000;
11113 : 00000;
11114 : 00000;
11115 : 00000;
11116 : 00000;
11117 : 00000;
11120 : 00000;
11121 : 00000;
11122 : 00000;
11123 : 00000;
11124 : 00000;
11125 : 00000;
11126 : 00000;
11127 : 00000;
11130 : 00000;
11131 : 00000;
11132 : 00000;
11133 : 00000;
11134 : 00000;
11135 : 00000;
11136 : 00000;
11137 : 00000;
11140 : 00000;
11141 : 00000;
11142 : 00000;
11143 : 00000;
11144 : 00000;
11145 : 00000;
11146 : 00000;
11147 : 00000;
11150 : 00000;
11151 : 00000;
11152 : 00000;
11153 : 00000;
11154 : 00000;
11155 : 00000;
11156 : 00000;
11157 : 00000;
11160 : 00000;
11161 : 00000;
11162 : 00000;
11163 : 00000;
11164 : 00000;
11165 : 00000;
11166 : 00000;
11167 : 00000;
11170 : 00000;
11171 : 00000;
11172 : 00000;
11173 : 00000;
11174 : 00000;
11175 : 00000;
11176 : 00000;
11177 : 00000;
11200 : 00000;
11201 : 00000;
11202 : 00000;
11203 : 00000;
11204 : 00000;
11205 : 00000;
11206 : 00000;
11207 : 00000;
11210 : 00000;
11211 : 00000;
11212 : 00000;
11213 : 00000;
11214 : 00000;
11215 : 00000;
11216 : 00000;
11217 : 00000;
11220 : 00000;
11221 : 00000;
11222 : 00000;
11223 : 00000;
11224 : 00000;
11225 : 00000;
11226 : 00000;
11227 : 00000;
11230 : 00000;
11231 : 00000;
11232 : 00000;
11233 : 00000;
11234 : 00000;
11235 : 00000;
11236 : 00000;
11237 : 00000;
11240 : 00000;
11241 : 00000;
11242 : 00000;
11243 : 00000;
11244 : 00000;
11245 : 00000;
11246 : 00000;
11247 : 00000;
11250 : 00000;
11251 : 00000;
11252 : 00000;
11253 : 00000;
11254 : 00000;
11255 : 00000;
11256 : 00000;
11257 : 00000;
11260 : 00000;
11261 : 00000;
11262 : 00000;
11263 : 00000;
11264 : 00000;
11265 : 00000;
11266 : 00000;
11267 : 00000;
11270 : 00000;
11271 : 00000;
11272 : 00000;
11273 : 00000;
11274 : 00000;
11275 : 00000;
11276 : 00000;
11277 : 00000;
11300 : 00000;
11301 : 00000;
11302 : 00000;
11303 : 00000;
11304 : 00000;
11305 : 00000;
11306 : 00000;
11307 : 00000;
11310 : 00000;
11311 : 00000;
11312 : 00000;
11313 : 00000;
11314 : 00000;
11315 : 00000;
11316 : 00000;
11317 : 00000;
11320 : 00000;
11321 : 00000;
11322 : 00000;
11323 : 00000;
11324 : 00000;
11325 : 00000;
11326 : 00000;
11327 : 00000;
11330 : 00000;
11331 : 00000;
11332 : 00000;
11333 : 00000;
11334 : 00000;
11335 : 00000;
11336 : 00000;
11337 : 00000;
11340 : 00000;
11341 : 00000;
11342 : 00000;
11343 : 00000;
11344 : 00000;
11345 : 00000;
11346 : 00000;
11347 : 00000;
11350 : 00000;
11351 : 00000;
11352 : 00000;
11353 : 00000;
11354 : 00000;
11355 : 00000;
11356 : 00000;
11357 : 00000;
11360 : 00000;
11361 : 00000;
11362 : 00000;
11363 : 00000;
11364 : 00000;
11365 : 00000;
11366 : 00000;
11367 : 00000;
11370 : 00000;
11371 : 00000;
11372 : 00000;
11373 : 00000;
11374 : 00000;
11375 : 00000;
11376 : 00000;
11377 : 00000;
11400 : 00000;
11401 : 00000;
11402 : 00000;
11403 : 00000;
11404 : 00000;
11405 : 00000;
11406 : 00000;
11407 : 00000;
11410 : 00000;
11411 : 00000;
11412 : 00000;
11413 : 00000;
11414 : 00000;
11415 : 00000;
11416 : 00000;
11417 : 00000;
11420 : 00000;
11421 : 00000;
11422 : 00000;
11423 : 00000;
11424 : 00000;
11425 : 00000;
11426 : 00000;
11427 : 00000;
11430 : 00000;
11431 : 00000;
11432 : 00000;
11433 : 00000;
11434 : 00000;
11435 : 00000;
11436 : 00000;
11437 : 00000;
11440 : 00000;
11441 : 00000;
11442 : 00000;
11443 : 00000;
11444 : 00000;
11445 : 00000;
11446 : 00000;
11447 : 00000;
11450 : 00000;
11451 : 00000;
11452 : 00000;
11453 : 00000;
11454 : 00000;
11455 : 00000;
11456 : 00000;
11457 : 00000;
11460 : 00000;
11461 : 00000;
11462 : 00000;
11463 : 00000;
11464 : 00000;
11465 : 00000;
11466 : 00000;
11467 : 00000;
11470 : 00000;
11471 : 00000;
11472 : 00000;
11473 : 00000;
11474 : 00000;
11475 : 00000;
11476 : 00000;
11477 : 00000;
11500 : 00000;
11501 : 00000;
11502 : 00000;
11503 : 00000;
11504 : 00000;
11505 : 00000;
11506 : 00000;
11507 : 00000;
11510 : 00000;
11511 : 00000;
11512 : 00000;
11513 : 00000;
11514 : 00000;
11515 : 00000;
11516 : 00000;
11517 : 00000;
11520 : 00000;
11521 : 00000;
11522 : 00000;
11523 : 00000;
11524 : 00000;
11525 : 00000;
11526 : 00000;
11527 : 00000;
11530 : 00000;
11531 : 00000;
11532 : 00000;
11533 : 00000;
11534 : 00000;
11535 : 00000;
11536 : 00000;
11537 : 00000;
11540 : 00000;
11541 : 00000;
11542 : 00000;
11543 : 00000;
11544 : 00000;
11545 : 00000;
11546 : 00000;
11547 : 00000;
11550 : 00000;
11551 : 00000;
11552 : 00000;
11553 : 00000;
11554 : 00000;
11555 : 00000;
11556 : 00000;
11557 : 00000;
11560 : 00000;
11561 : 00000;
11562 : 00000;
11563 : 00000;
11564 : 00000;
11565 : 00000;
11566 : 00000;
11567 : 00000;
11570 : 00000;
11571 : 00000;
11572 : 00000;
11573 : 00000;
11574 : 00000;
11575 : 00000;
11576 : 00000;
11577 : 00000;
11600 : 00000;
11601 : 00000;
11602 : 00000;
11603 : 00000;
11604 : 00000;
11605 : 00000;
11606 : 00000;
11607 : 00000;
11610 : 00000;
11611 : 00000;
11612 : 00000;
11613 : 00000;
11614 : 00000;
11615 : 00000;
11616 : 00000;
11617 : 00000;
11620 : 00000;
11621 : 00000;
11622 : 00000;
11623 : 00000;
11624 : 00000;
11625 : 00000;
11626 : 00000;
11627 : 00000;
11630 : 00000;
11631 : 00000;
11632 : 00000;
11633 : 00000;
11634 : 00000;
11635 : 00000;
11636 : 00000;
11637 : 00000;
11640 : 00000;
11641 : 00000;
11642 : 00000;
11643 : 00000;
11644 : 00000;
11645 : 00000;
11646 : 00000;
11647 : 00000;
11650 : 00000;
11651 : 00000;
11652 : 00000;
11653 : 00000;
11654 : 00000;
11655 : 00000;
11656 : 00000;
11657 : 00000;
11660 : 00000;
11661 : 00000;
11662 : 00000;
11663 : 00000;
11664 : 00000;
11665 : 00000;
11666 : 00000;
11667 : 00000;
11670 : 00000;
11671 : 00000;
11672 : 00000;
11673 : 00000;
11674 : 00000;
11675 : 00000;
11676 : 00000;
11677 : 00000;
11700 : 00000;
11701 : 00000;
11702 : 00000;
11703 : 00000;
11704 : 00000;
11705 : 00000;
11706 : 00000;
11707 : 00000;
11710 : 00000;
11711 : 00000;
11712 : 00000;
11713 : 00000;
11714 : 00000;
11715 : 00000;
11716 : 00000;
11717 : 00000;
11720 : 00000;
11721 : 00000;
11722 : 00000;
11723 : 00000;
11724 : 00000;
11725 : 00000;
11726 : 00000;
11727 : 00000;
11730 : 00000;
11731 : 00000;
11732 : 00000;
11733 : 00000;
11734 : 00000;
11735 : 00000;
11736 : 00000;
11737 : 00000;
11740 : 00000;
11741 : 00000;
11742 : 00000;
11743 : 00000;
11744 : 00000;
11745 : 00000;
11746 : 00000;
11747 : 00000;
11750 : 00000;
11751 : 00000;
11752 : 00000;
11753 : 00000;
11754 : 00000;
11755 : 00000;
11756 : 00000;
11757 : 00000;
11760 : 00000;
11761 : 00000;
11762 : 00000;
11763 : 00000;
11764 : 00000;
11765 : 00000;
11766 : 00000;
11767 : 00000;
11770 : 00000;
11771 : 00000;
11772 : 00000;
11773 : 00000;
11774 : 00000;
11775 : 00000;
11776 : 00000;
11777 : 00000;
12000 : 00000;
12001 : 00000;
12002 : 00000;
12003 : 00000;
12004 : 00000;
12005 : 00000;
12006 : 00000;
12007 : 00000;
12010 : 00000;
12011 : 00000;
12012 : 00000;
12013 : 00000;
12014 : 00000;
12015 : 00000;
12016 : 00000;
12017 : 00000;
12020 : 00000;
12021 : 00000;
12022 : 00000;
12023 : 00000;
12024 : 00000;
12025 : 00000;
12026 : 00000;
12027 : 00000;
12030 : 00000;
12031 : 00000;
12032 : 00000;
12033 : 00000;
12034 : 00000;
12035 : 00000;
12036 : 00000;
12037 : 00000;
12040 : 00000;
12041 : 00000;
12042 : 00000;
12043 : 00000;
12044 : 00000;
12045 : 00000;
12046 : 00000;
12047 : 00000;
12050 : 00000;
12051 : 00000;
12052 : 00000;
12053 : 00000;
12054 : 00000;
12055 : 00000;
12056 : 00000;
12057 : 00000;
12060 : 00000;
12061 : 00000;
12062 : 00000;
12063 : 00000;
12064 : 00000;
12065 : 00000;
12066 : 00000;
12067 : 00000;
12070 : 00000;
12071 : 00000;
12072 : 00000;
12073 : 00000;
12074 : 00000;
12075 : 00000;
12076 : 00000;
12077 : 00000;
12100 : 00000;
12101 : 00000;
12102 : 00000;
12103 : 00000;
12104 : 00000;
12105 : 00000;
12106 : 00000;
12107 : 00000;
12110 : 00000;
12111 : 00000;
12112 : 00000;
12113 : 00000;
12114 : 00000;
12115 : 00000;
12116 : 00000;
12117 : 00000;
12120 : 00000;
12121 : 00000;
12122 : 00000;
12123 : 00000;
12124 : 00000;
12125 : 00000;
12126 : 00000;
12127 : 00000;
12130 : 00000;
12131 : 00000;
12132 : 00000;
12133 : 00000;
12134 : 00000;
12135 : 00000;
12136 : 00000;
12137 : 00000;
12140 : 00000;
12141 : 00000;
12142 : 00000;
12143 : 00000;
12144 : 00000;
12145 : 00000;
12146 : 00000;
12147 : 00000;
12150 : 00000;
12151 : 00000;
12152 : 00000;
12153 : 00000;
12154 : 00000;
12155 : 00000;
12156 : 00000;
12157 : 00000;
12160 : 00000;
12161 : 00000;
12162 : 00000;
12163 : 00000;
12164 : 00000;
12165 : 00000;
12166 : 00000;
12167 : 00000;
12170 : 00000;
12171 : 00000;
12172 : 00000;
12173 : 00000;
12174 : 00000;
12175 : 00000;
12176 : 00000;
12177 : 00000;
12200 : 00000;
12201 : 00000;
12202 : 00000;
12203 : 00000;
12204 : 00000;
12205 : 00000;
12206 : 00000;
12207 : 00000;
12210 : 00000;
12211 : 00000;
12212 : 00000;
12213 : 00000;
12214 : 00000;
12215 : 00000;
12216 : 00000;
12217 : 00000;
12220 : 00000;
12221 : 00000;
12222 : 00000;
12223 : 00000;
12224 : 00000;
12225 : 00000;
12226 : 00000;
12227 : 00000;
12230 : 00000;
12231 : 00000;
12232 : 00000;
12233 : 00000;
12234 : 00000;
12235 : 00000;
12236 : 00000;
12237 : 00000;
12240 : 00000;
12241 : 00000;
12242 : 00000;
12243 : 00000;
12244 : 00000;
12245 : 00000;
12246 : 00000;
12247 : 00000;
12250 : 00000;
12251 : 00000;
12252 : 00000;
12253 : 00000;
12254 : 00000;
12255 : 00000;
12256 : 00000;
12257 : 00000;
12260 : 00000;
12261 : 00000;
12262 : 00000;
12263 : 00000;
12264 : 00000;
12265 : 00000;
12266 : 00000;
12267 : 00000;
12270 : 00000;
12271 : 00000;
12272 : 00000;
12273 : 00000;
12274 : 00000;
12275 : 00000;
12276 : 00000;
12277 : 00000;
12300 : 00000;
12301 : 00000;
12302 : 00000;
12303 : 00000;
12304 : 00000;
12305 : 00000;
12306 : 00000;
12307 : 00000;
12310 : 00000;
12311 : 00000;
12312 : 00000;
12313 : 00000;
12314 : 00000;
12315 : 00000;
12316 : 00000;
12317 : 00000;
12320 : 00000;
12321 : 00000;
12322 : 00000;
12323 : 00000;
12324 : 00000;
12325 : 00000;
12326 : 00000;
12327 : 00000;
12330 : 00000;
12331 : 00000;
12332 : 00000;
12333 : 00000;
12334 : 00000;
12335 : 00000;
12336 : 00000;
12337 : 00000;
12340 : 00000;
12341 : 00000;
12342 : 00000;
12343 : 00000;
12344 : 00000;
12345 : 00000;
12346 : 00000;
12347 : 00000;
12350 : 00000;
12351 : 00000;
12352 : 00000;
12353 : 00000;
12354 : 00000;
12355 : 00000;
12356 : 00000;
12357 : 00000;
12360 : 00000;
12361 : 00000;
12362 : 00000;
12363 : 00000;
12364 : 00000;
12365 : 00000;
12366 : 00000;
12367 : 00000;
12370 : 00000;
12371 : 00000;
12372 : 00000;
12373 : 00000;
12374 : 00000;
12375 : 00000;
12376 : 00000;
12377 : 00000;
12400 : 00000;
12401 : 00000;
12402 : 00000;
12403 : 00000;
12404 : 00000;
12405 : 00000;
12406 : 00000;
12407 : 00000;
12410 : 00000;
12411 : 00000;
12412 : 00000;
12413 : 00000;
12414 : 00000;
12415 : 00000;
12416 : 00000;
12417 : 00000;
12420 : 00000;
12421 : 00000;
12422 : 00000;
12423 : 00000;
12424 : 00000;
12425 : 00000;
12426 : 00000;
12427 : 00000;
12430 : 00000;
12431 : 00000;
12432 : 00000;
12433 : 00000;
12434 : 00000;
12435 : 00000;
12436 : 00000;
12437 : 00000;
12440 : 00000;
12441 : 00000;
12442 : 00000;
12443 : 00000;
12444 : 00000;
12445 : 00000;
12446 : 00000;
12447 : 00000;
12450 : 00000;
12451 : 00000;
12452 : 00000;
12453 : 00000;
12454 : 00000;
12455 : 00000;
12456 : 00000;
12457 : 00000;
12460 : 00000;
12461 : 00000;
12462 : 00000;
12463 : 00000;
12464 : 00000;
12465 : 00000;
12466 : 00000;
12467 : 00000;
12470 : 00000;
12471 : 00000;
12472 : 00000;
12473 : 00000;
12474 : 00000;
12475 : 00000;
12476 : 00000;
12477 : 00000;
12500 : 00000;
12501 : 00000;
12502 : 00000;
12503 : 00000;
12504 : 00000;
12505 : 00000;
12506 : 00000;
12507 : 00000;
12510 : 00000;
12511 : 00000;
12512 : 00000;
12513 : 00000;
12514 : 00000;
12515 : 00000;
12516 : 00000;
12517 : 00000;
12520 : 00000;
12521 : 00000;
12522 : 00000;
12523 : 00000;
12524 : 00000;
12525 : 00000;
12526 : 00000;
12527 : 00000;
12530 : 00000;
12531 : 00000;
12532 : 00000;
12533 : 00000;
12534 : 00000;
12535 : 00000;
12536 : 00000;
12537 : 00000;
12540 : 00000;
12541 : 00000;
12542 : 00000;
12543 : 00000;
12544 : 00000;
12545 : 00000;
12546 : 00000;
12547 : 00000;
12550 : 00000;
12551 : 00000;
12552 : 00000;
12553 : 00000;
12554 : 00000;
12555 : 00000;
12556 : 00000;
12557 : 00000;
12560 : 00000;
12561 : 00000;
12562 : 00000;
12563 : 00000;
12564 : 00000;
12565 : 00000;
12566 : 00000;
12567 : 00000;
12570 : 00000;
12571 : 00000;
12572 : 00000;
12573 : 00000;
12574 : 00000;
12575 : 00000;
12576 : 00000;
12577 : 00000;
12600 : 00000;
12601 : 00000;
12602 : 00000;
12603 : 00000;
12604 : 00000;
12605 : 00000;
12606 : 00000;
12607 : 00000;
12610 : 00000;
12611 : 00000;
12612 : 00000;
12613 : 00000;
12614 : 00000;
12615 : 00000;
12616 : 00000;
12617 : 00000;
12620 : 00000;
12621 : 00000;
12622 : 00000;
12623 : 00000;
12624 : 00000;
12625 : 00000;
12626 : 00000;
12627 : 00000;
12630 : 00000;
12631 : 00000;
12632 : 00000;
12633 : 00000;
12634 : 00000;
12635 : 00000;
12636 : 00000;
12637 : 00000;
12640 : 00000;
12641 : 00000;
12642 : 00000;
12643 : 00000;
12644 : 00000;
12645 : 00000;
12646 : 00000;
12647 : 00000;
12650 : 00000;
12651 : 00000;
12652 : 00000;
12653 : 00000;
12654 : 00000;
12655 : 00000;
12656 : 00000;
12657 : 00000;
12660 : 00000;
12661 : 00000;
12662 : 00000;
12663 : 00000;
12664 : 00000;
12665 : 00000;
12666 : 00000;
12667 : 00000;
12670 : 00000;
12671 : 00000;
12672 : 00000;
12673 : 00000;
12674 : 00000;
12675 : 00000;
12676 : 00000;
12677 : 00000;
12700 : 00000;
12701 : 00000;
12702 : 00000;
12703 : 00000;
12704 : 00000;
12705 : 00000;
12706 : 00000;
12707 : 00000;
12710 : 00000;
12711 : 00000;
12712 : 00000;
12713 : 00000;
12714 : 00000;
12715 : 00000;
12716 : 00000;
12717 : 00000;
12720 : 00000;
12721 : 00000;
12722 : 00000;
12723 : 00000;
12724 : 00000;
12725 : 00000;
12726 : 00000;
12727 : 00000;
12730 : 00000;
12731 : 00000;
12732 : 00000;
12733 : 00000;
12734 : 00000;
12735 : 00000;
12736 : 00000;
12737 : 00000;
12740 : 00000;
12741 : 00000;
12742 : 00000;
12743 : 00000;
12744 : 00000;
12745 : 00000;
12746 : 00000;
12747 : 00000;
12750 : 00000;
12751 : 00000;
12752 : 00000;
12753 : 00000;
12754 : 00000;
12755 : 00000;
12756 : 00000;
12757 : 00000;
12760 : 00000;
12761 : 00000;
12762 : 00000;
12763 : 00000;
12764 : 00000;
12765 : 00000;
12766 : 00000;
12767 : 00000;
12770 : 00000;
12771 : 00000;
12772 : 00000;
12773 : 00000;
12774 : 00000;
12775 : 00000;
12776 : 00000;
12777 : 00000;
13000 : 00000;
13001 : 00000;
13002 : 00000;
13003 : 00000;
13004 : 00000;
13005 : 00000;
13006 : 00000;
13007 : 00000;
13010 : 00000;
13011 : 00000;
13012 : 00000;
13013 : 00000;
13014 : 00000;
13015 : 00000;
13016 : 00000;
13017 : 00000;
13020 : 00000;
13021 : 00000;
13022 : 00000;
13023 : 00000;
13024 : 00000;
13025 : 00000;
13026 : 00000;
13027 : 00000;
13030 : 00000;
13031 : 00000;
13032 : 00000;
13033 : 00000;
13034 : 00000;
13035 : 00000;
13036 : 00000;
13037 : 00000;
13040 : 00000;
13041 : 00000;
13042 : 00000;
13043 : 00000;
13044 : 00000;
13045 : 00000;
13046 : 00000;
13047 : 00000;
13050 : 00000;
13051 : 00000;
13052 : 00000;
13053 : 00000;
13054 : 00000;
13055 : 00000;
13056 : 00000;
13057 : 00000;
13060 : 00000;
13061 : 00000;
13062 : 00000;
13063 : 00000;
13064 : 00000;
13065 : 00000;
13066 : 00000;
13067 : 00000;
13070 : 00000;
13071 : 00000;
13072 : 00000;
13073 : 00000;
13074 : 00000;
13075 : 00000;
13076 : 00000;
13077 : 00000;
13100 : 00000;
13101 : 00000;
13102 : 00000;
13103 : 00000;
13104 : 00000;
13105 : 00000;
13106 : 00000;
13107 : 00000;
13110 : 00000;
13111 : 00000;
13112 : 00000;
13113 : 00000;
13114 : 00000;
13115 : 00000;
13116 : 00000;
13117 : 00000;
13120 : 00000;
13121 : 00000;
13122 : 00000;
13123 : 00000;
13124 : 00000;
13125 : 00000;
13126 : 00000;
13127 : 00000;
13130 : 00000;
13131 : 00000;
13132 : 00000;
13133 : 00000;
13134 : 00000;
13135 : 00000;
13136 : 00000;
13137 : 00000;
13140 : 00000;
13141 : 00000;
13142 : 00000;
13143 : 00000;
13144 : 00000;
13145 : 00000;
13146 : 00000;
13147 : 00000;
13150 : 00000;
13151 : 00000;
13152 : 00000;
13153 : 00000;
13154 : 00000;
13155 : 00000;
13156 : 00000;
13157 : 00000;
13160 : 00000;
13161 : 00000;
13162 : 00000;
13163 : 00000;
13164 : 00000;
13165 : 00000;
13166 : 00000;
13167 : 00000;
13170 : 00000;
13171 : 00000;
13172 : 00000;
13173 : 00000;
13174 : 00000;
13175 : 00000;
13176 : 00000;
13177 : 00000;
13200 : 00000;
13201 : 00000;
13202 : 00000;
13203 : 00000;
13204 : 00000;
13205 : 00000;
13206 : 00000;
13207 : 00000;
13210 : 00000;
13211 : 00000;
13212 : 00000;
13213 : 00000;
13214 : 00000;
13215 : 00000;
13216 : 00000;
13217 : 00000;
13220 : 00000;
13221 : 00000;
13222 : 00000;
13223 : 00000;
13224 : 00000;
13225 : 00000;
13226 : 00000;
13227 : 00000;
13230 : 00000;
13231 : 00000;
13232 : 00000;
13233 : 00000;
13234 : 00000;
13235 : 00000;
13236 : 00000;
13237 : 00000;
13240 : 00000;
13241 : 00000;
13242 : 00000;
13243 : 00000;
13244 : 00000;
13245 : 00000;
13246 : 00000;
13247 : 00000;
13250 : 00000;
13251 : 00000;
13252 : 00000;
13253 : 00000;
13254 : 00000;
13255 : 00000;
13256 : 00000;
13257 : 00000;
13260 : 00000;
13261 : 00000;
13262 : 00000;
13263 : 00000;
13264 : 00000;
13265 : 00000;
13266 : 00000;
13267 : 00000;
13270 : 00000;
13271 : 00000;
13272 : 00000;
13273 : 00000;
13274 : 00000;
13275 : 00000;
13276 : 00000;
13277 : 00000;
13300 : 00000;
13301 : 00000;
13302 : 00000;
13303 : 00000;
13304 : 00000;
13305 : 00000;
13306 : 00000;
13307 : 00000;
13310 : 00000;
13311 : 00000;
13312 : 00000;
13313 : 00000;
13314 : 00000;
13315 : 00000;
13316 : 00000;
13317 : 00000;
13320 : 00000;
13321 : 00000;
13322 : 00000;
13323 : 00000;
13324 : 00000;
13325 : 00000;
13326 : 00000;
13327 : 00000;
13330 : 00000;
13331 : 00000;
13332 : 00000;
13333 : 00000;
13334 : 00000;
13335 : 00000;
13336 : 00000;
13337 : 00000;
13340 : 00000;
13341 : 00000;
13342 : 00000;
13343 : 00000;
13344 : 00000;
13345 : 00000;
13346 : 00000;
13347 : 00000;
13350 : 00000;
13351 : 00000;
13352 : 00000;
13353 : 00000;
13354 : 00000;
13355 : 00000;
13356 : 00000;
13357 : 00000;
13360 : 00000;
13361 : 00000;
13362 : 00000;
13363 : 00000;
13364 : 00000;
13365 : 00000;
13366 : 00000;
13367 : 00000;
13370 : 00000;
13371 : 00000;
13372 : 00000;
13373 : 00000;
13374 : 00000;
13375 : 00000;
13376 : 00000;
13377 : 00000;
13400 : 00000;
13401 : 00000;
13402 : 00000;
13403 : 00000;
13404 : 00000;
13405 : 00000;
13406 : 00000;
13407 : 00000;
13410 : 00000;
13411 : 00000;
13412 : 00000;
13413 : 00000;
13414 : 00000;
13415 : 00000;
13416 : 00000;
13417 : 00000;
13420 : 00000;
13421 : 00000;
13422 : 00000;
13423 : 00000;
13424 : 00000;
13425 : 00000;
13426 : 00000;
13427 : 00000;
13430 : 00000;
13431 : 00000;
13432 : 00000;
13433 : 00000;
13434 : 00000;
13435 : 00000;
13436 : 00000;
13437 : 00000;
13440 : 00000;
13441 : 00000;
13442 : 00000;
13443 : 00000;
13444 : 00000;
13445 : 00000;
13446 : 00000;
13447 : 00000;
13450 : 00000;
13451 : 00000;
13452 : 00000;
13453 : 00000;
13454 : 00000;
13455 : 00000;
13456 : 00000;
13457 : 00000;
13460 : 00000;
13461 : 00000;
13462 : 00000;
13463 : 00000;
13464 : 00000;
13465 : 00000;
13466 : 00000;
13467 : 00000;
13470 : 00000;
13471 : 00000;
13472 : 00000;
13473 : 00000;
13474 : 00000;
13475 : 00000;
13476 : 00000;
13477 : 00000;
13500 : 00000;
13501 : 00000;
13502 : 00000;
13503 : 00000;
13504 : 00000;
13505 : 00000;
13506 : 00000;
13507 : 00000;
13510 : 00000;
13511 : 00000;
13512 : 00000;
13513 : 00000;
13514 : 00000;
13515 : 00000;
13516 : 00000;
13517 : 00000;
13520 : 00000;
13521 : 00000;
13522 : 00000;
13523 : 00000;
13524 : 00000;
13525 : 00000;
13526 : 00000;
13527 : 00000;
13530 : 00000;
13531 : 00000;
13532 : 00000;
13533 : 00000;
13534 : 00000;
13535 : 00000;
13536 : 00000;
13537 : 00000;
13540 : 00000;
13541 : 00000;
13542 : 00000;
13543 : 00000;
13544 : 00000;
13545 : 00000;
13546 : 00000;
13547 : 00000;
13550 : 00000;
13551 : 00000;
13552 : 00000;
13553 : 00000;
13554 : 00000;
13555 : 00000;
13556 : 00000;
13557 : 00000;
13560 : 00000;
13561 : 00000;
13562 : 00000;
13563 : 00000;
13564 : 00000;
13565 : 00000;
13566 : 00000;
13567 : 00000;
13570 : 00000;
13571 : 00000;
13572 : 00000;
13573 : 00000;
13574 : 00000;
13575 : 00000;
13576 : 00000;
13577 : 00000;
13600 : 00000;
13601 : 00000;
13602 : 00000;
13603 : 00000;
13604 : 00000;
13605 : 00000;
13606 : 00000;
13607 : 00000;
13610 : 00000;
13611 : 00000;
13612 : 00000;
13613 : 00000;
13614 : 00000;
13615 : 00000;
13616 : 00000;
13617 : 00000;
13620 : 00000;
13621 : 00000;
13622 : 00000;
13623 : 00000;
13624 : 00000;
13625 : 00000;
13626 : 00000;
13627 : 00000;
13630 : 00000;
13631 : 00000;
13632 : 00000;
13633 : 00000;
13634 : 00000;
13635 : 00000;
13636 : 00000;
13637 : 00000;
13640 : 00000;
13641 : 00000;
13642 : 00000;
13643 : 00000;
13644 : 00000;
13645 : 00000;
13646 : 00000;
13647 : 00000;
13650 : 00000;
13651 : 00000;
13652 : 00000;
13653 : 00000;
13654 : 00000;
13655 : 00000;
13656 : 00000;
13657 : 00000;
13660 : 00000;
13661 : 00000;
13662 : 00000;
13663 : 00000;
13664 : 00000;
13665 : 00000;
13666 : 00000;
13667 : 00000;
13670 : 00000;
13671 : 00000;
13672 : 00000;
13673 : 00000;
13674 : 00000;
13675 : 00000;
13676 : 00000;
13677 : 00000;
13700 : 00000;
13701 : 00000;
13702 : 00000;
13703 : 00000;
13704 : 00000;
13705 : 00000;
13706 : 00000;
13707 : 00000;
13710 : 00000;
13711 : 00000;
13712 : 00000;
13713 : 00000;
13714 : 00000;
13715 : 00000;
13716 : 00000;
13717 : 00000;
13720 : 00000;
13721 : 00000;
13722 : 00000;
13723 : 00000;
13724 : 00000;
13725 : 00000;
13726 : 00000;
13727 : 00000;
13730 : 00000;
13731 : 00000;
13732 : 00000;
13733 : 00000;
13734 : 00000;
13735 : 00000;
13736 : 00000;
13737 : 00000;
13740 : 00000;
13741 : 00000;
13742 : 00000;
13743 : 00000;
13744 : 00000;
13745 : 00000;
13746 : 00000;
13747 : 00000;
13750 : 00000;
13751 : 00000;
13752 : 00000;
13753 : 00000;
13754 : 00000;
13755 : 00000;
13756 : 00000;
13757 : 00000;
13760 : 00000;
13761 : 00000;
13762 : 00000;
13763 : 00000;
13764 : 00000;
13765 : 00000;
13766 : 00000;
13767 : 00000;
13770 : 00000;
13771 : 00000;
13772 : 00000;
13773 : 00000;
13774 : 00000;
13775 : 00000;
13776 : 00000;
13777 : 00000;
14000 : 00000;
14001 : 00000;
14002 : 00000;
14003 : 00000;
14004 : 00000;
14005 : 00000;
14006 : 00000;
14007 : 00000;
14010 : 00000;
14011 : 00000;
14012 : 00000;
14013 : 00000;
14014 : 00000;
14015 : 00000;
14016 : 00000;
14017 : 00000;
14020 : 00000;
14021 : 00000;
14022 : 00000;
14023 : 00000;
14024 : 00000;
14025 : 00000;
14026 : 00000;
14027 : 00000;
14030 : 00000;
14031 : 00000;
14032 : 00000;
14033 : 00000;
14034 : 00000;
14035 : 00000;
14036 : 00000;
14037 : 00000;
14040 : 00000;
14041 : 00000;
14042 : 00000;
14043 : 00000;
14044 : 00000;
14045 : 00000;
14046 : 00000;
14047 : 00000;
14050 : 00000;
14051 : 00000;
14052 : 00000;
14053 : 00000;
14054 : 00000;
14055 : 00000;
14056 : 00000;
14057 : 00000;
14060 : 00000;
14061 : 00000;
14062 : 00000;
14063 : 00000;
14064 : 00000;
14065 : 00000;
14066 : 00000;
14067 : 00000;
14070 : 00000;
14071 : 00000;
14072 : 00000;
14073 : 00000;
14074 : 00000;
14075 : 00000;
14076 : 00000;
14077 : 00000;
14100 : 00000;
14101 : 00000;
14102 : 00000;
14103 : 00000;
14104 : 00000;
14105 : 00000;
14106 : 00000;
14107 : 00000;
14110 : 00000;
14111 : 00000;
14112 : 00000;
14113 : 00000;
14114 : 00000;
14115 : 00000;
14116 : 00000;
14117 : 00000;
14120 : 00000;
14121 : 00000;
14122 : 00000;
14123 : 00000;
14124 : 00000;
14125 : 00000;
14126 : 00000;
14127 : 00000;
14130 : 00000;
14131 : 00000;
14132 : 00000;
14133 : 00000;
14134 : 00000;
14135 : 00000;
14136 : 00000;
14137 : 00000;
14140 : 00000;
14141 : 00000;
14142 : 00000;
14143 : 00000;
14144 : 00000;
14145 : 00000;
14146 : 00000;
14147 : 00000;
14150 : 00000;
14151 : 00000;
14152 : 00000;
14153 : 00000;
14154 : 00000;
14155 : 00000;
14156 : 00000;
14157 : 00000;
14160 : 00000;
14161 : 00000;
14162 : 00000;
14163 : 00000;
14164 : 00000;
14165 : 00000;
14166 : 00000;
14167 : 00000;
14170 : 00000;
14171 : 00000;
14172 : 00000;
14173 : 00000;
14174 : 00000;
14175 : 00000;
14176 : 00000;
14177 : 00000;
14200 : 00000;
14201 : 00000;
14202 : 00000;
14203 : 00000;
14204 : 00000;
14205 : 00000;
14206 : 00000;
14207 : 00000;
14210 : 00000;
14211 : 00000;
14212 : 00000;
14213 : 00000;
14214 : 00000;
14215 : 00000;
14216 : 00000;
14217 : 00000;
14220 : 00000;
14221 : 00000;
14222 : 00000;
14223 : 00000;
14224 : 00000;
14225 : 00000;
14226 : 00000;
14227 : 00000;
14230 : 00000;
14231 : 00000;
14232 : 00000;
14233 : 00000;
14234 : 00000;
14235 : 00000;
14236 : 00000;
14237 : 00000;
14240 : 00000;
14241 : 00000;
14242 : 00000;
14243 : 00000;
14244 : 00000;
14245 : 00000;
14246 : 00000;
14247 : 00000;
14250 : 00000;
14251 : 00000;
14252 : 00000;
14253 : 00000;
14254 : 00000;
14255 : 00000;
14256 : 00000;
14257 : 00000;
14260 : 00000;
14261 : 00000;
14262 : 00000;
14263 : 00000;
14264 : 00000;
14265 : 00000;
14266 : 00000;
14267 : 00000;
14270 : 00000;
14271 : 00000;
14272 : 00000;
14273 : 00000;
14274 : 00000;
14275 : 00000;
14276 : 00000;
14277 : 00000;
14300 : 00000;
14301 : 00000;
14302 : 00000;
14303 : 00000;
14304 : 00000;
14305 : 00000;
14306 : 00000;
14307 : 00000;
14310 : 00000;
14311 : 00000;
14312 : 00000;
14313 : 00000;
14314 : 00000;
14315 : 00000;
14316 : 00000;
14317 : 00000;
14320 : 00000;
14321 : 00000;
14322 : 00000;
14323 : 00000;
14324 : 00000;
14325 : 00000;
14326 : 00000;
14327 : 00000;
14330 : 00000;
14331 : 00000;
14332 : 00000;
14333 : 00000;
14334 : 00000;
14335 : 00000;
14336 : 00000;
14337 : 00000;
14340 : 00000;
14341 : 00000;
14342 : 00000;
14343 : 00000;
14344 : 00000;
14345 : 00000;
14346 : 00000;
14347 : 00000;
14350 : 00000;
14351 : 00000;
14352 : 00000;
14353 : 00000;
14354 : 00000;
14355 : 00000;
14356 : 00000;
14357 : 00000;
14360 : 00000;
14361 : 00000;
14362 : 00000;
14363 : 00000;
14364 : 00000;
14365 : 00000;
14366 : 00000;
14367 : 00000;
14370 : 00000;
14371 : 00000;
14372 : 00000;
14373 : 00000;
14374 : 00000;
14375 : 00000;
14376 : 00000;
14377 : 00000;
14400 : 00000;
14401 : 00000;
14402 : 00000;
14403 : 00000;
14404 : 00000;
14405 : 00000;
14406 : 00000;
14407 : 00000;
14410 : 00000;
14411 : 00000;
14412 : 00000;
14413 : 00000;
14414 : 00000;
14415 : 00000;
14416 : 00000;
14417 : 00000;
14420 : 00000;
14421 : 00000;
14422 : 00000;
14423 : 00000;
14424 : 00000;
14425 : 00000;
14426 : 00000;
14427 : 00000;
14430 : 00000;
14431 : 00000;
14432 : 00000;
14433 : 00000;
14434 : 00000;
14435 : 00000;
14436 : 00000;
14437 : 00000;
14440 : 00000;
14441 : 00000;
14442 : 00000;
14443 : 00000;
14444 : 00000;
14445 : 00000;
14446 : 00000;
14447 : 00000;
14450 : 00000;
14451 : 00000;
14452 : 00000;
14453 : 00000;
14454 : 00000;
14455 : 00000;
14456 : 00000;
14457 : 00000;
14460 : 00000;
14461 : 00000;
14462 : 00000;
14463 : 00000;
14464 : 00000;
14465 : 00000;
14466 : 00000;
14467 : 00000;
14470 : 00000;
14471 : 00000;
14472 : 00000;
14473 : 00000;
14474 : 00000;
14475 : 00000;
14476 : 00000;
14477 : 00000;
14500 : 00000;
14501 : 00000;
14502 : 00000;
14503 : 00000;
14504 : 00000;
14505 : 00000;
14506 : 00000;
14507 : 00000;
14510 : 00000;
14511 : 00000;
14512 : 00000;
14513 : 00000;
14514 : 00000;
14515 : 00000;
14516 : 00000;
14517 : 00000;
14520 : 00000;
14521 : 00000;
14522 : 00000;
14523 : 00000;
14524 : 00000;
14525 : 00000;
14526 : 00000;
14527 : 00000;
14530 : 00000;
14531 : 00000;
14532 : 00000;
14533 : 00000;
14534 : 00000;
14535 : 00000;
14536 : 00000;
14537 : 00000;
14540 : 00000;
14541 : 00000;
14542 : 00000;
14543 : 00000;
14544 : 00000;
14545 : 00000;
14546 : 00000;
14547 : 00000;
14550 : 00000;
14551 : 00000;
14552 : 00000;
14553 : 00000;
14554 : 00000;
14555 : 00000;
14556 : 00000;
14557 : 00000;
14560 : 00000;
14561 : 00000;
14562 : 00000;
14563 : 00000;
14564 : 00000;
14565 : 00000;
14566 : 00000;
14567 : 00000;
14570 : 00000;
14571 : 00000;
14572 : 00000;
14573 : 00000;
14574 : 00000;
14575 : 00000;
14576 : 00000;
14577 : 00000;
14600 : 00000;
14601 : 00000;
14602 : 00000;
14603 : 00000;
14604 : 00000;
14605 : 00000;
14606 : 00000;
14607 : 00000;
14610 : 00000;
14611 : 00000;
14612 : 00000;
14613 : 00000;
14614 : 00000;
14615 : 00000;
14616 : 00000;
14617 : 00000;
14620 : 00000;
14621 : 00000;
14622 : 00000;
14623 : 00000;
14624 : 00000;
14625 : 00000;
14626 : 00000;
14627 : 00000;
14630 : 00000;
14631 : 00000;
14632 : 00000;
14633 : 00000;
14634 : 00000;
14635 : 00000;
14636 : 00000;
14637 : 00000;
14640 : 00000;
14641 : 00000;
14642 : 00000;
14643 : 00000;
14644 : 00000;
14645 : 00000;
14646 : 00000;
14647 : 00000;
14650 : 00000;
14651 : 00000;
14652 : 00000;
14653 : 00000;
14654 : 00000;
14655 : 00000;
14656 : 00000;
14657 : 00000;
14660 : 00000;
14661 : 00000;
14662 : 00000;
14663 : 00000;
14664 : 00000;
14665 : 00000;
14666 : 00000;
14667 : 00000;
14670 : 00000;
14671 : 00000;
14672 : 00000;
14673 : 00000;
14674 : 00000;
14675 : 00000;
14676 : 00000;
14677 : 00000;
14700 : 00000;
14701 : 00000;
14702 : 00000;
14703 : 00000;
14704 : 00000;
14705 : 00000;
14706 : 00000;
14707 : 00000;
14710 : 00000;
14711 : 00000;
14712 : 00000;
14713 : 00000;
14714 : 00000;
14715 : 00000;
14716 : 00000;
14717 : 00000;
14720 : 00000;
14721 : 00000;
14722 : 00000;
14723 : 00000;
14724 : 00000;
14725 : 00000;
14726 : 00000;
14727 : 00000;
14730 : 00000;
14731 : 00000;
14732 : 00000;
14733 : 00000;
14734 : 00000;
14735 : 00000;
14736 : 00000;
14737 : 00000;
14740 : 00000;
14741 : 00000;
14742 : 00000;
14743 : 00000;
14744 : 00000;
14745 : 00000;
14746 : 00000;
14747 : 00000;
14750 : 00000;
14751 : 00000;
14752 : 00000;
14753 : 00000;
14754 : 00000;
14755 : 00000;
14756 : 00000;
14757 : 00000;
14760 : 00000;
14761 : 00000;
14762 : 00000;
14763 : 00000;
14764 : 00000;
14765 : 00000;
14766 : 00000;
14767 : 00000;
14770 : 00000;
14771 : 00000;
14772 : 00000;
14773 : 00000;
14774 : 00000;
14775 : 00000;
14776 : 00000;
14777 : 00000;
15000 : 00000;
15001 : 00000;
15002 : 00000;
15003 : 00000;
15004 : 00000;
15005 : 00000;
15006 : 00000;
15007 : 00000;
15010 : 00000;
15011 : 00000;
15012 : 00000;
15013 : 00000;
15014 : 00000;
15015 : 00000;
15016 : 00000;
15017 : 00000;
15020 : 00000;
15021 : 00000;
15022 : 00000;
15023 : 00000;
15024 : 00000;
15025 : 00000;
15026 : 00000;
15027 : 00000;
15030 : 00000;
15031 : 00000;
15032 : 00000;
15033 : 00000;
15034 : 00000;
15035 : 00000;
15036 : 00000;
15037 : 00000;
15040 : 00000;
15041 : 00000;
15042 : 00000;
15043 : 00000;
15044 : 00000;
15045 : 00000;
15046 : 00000;
15047 : 00000;
15050 : 00000;
15051 : 00000;
15052 : 00000;
15053 : 00000;
15054 : 00000;
15055 : 00000;
15056 : 00000;
15057 : 00000;
15060 : 00000;
15061 : 00000;
15062 : 00000;
15063 : 00000;
15064 : 00000;
15065 : 00000;
15066 : 00000;
15067 : 00000;
15070 : 00000;
15071 : 00000;
15072 : 00000;
15073 : 00000;
15074 : 00000;
15075 : 00000;
15076 : 00000;
15077 : 00000;
15100 : 00000;
15101 : 00000;
15102 : 00000;
15103 : 00000;
15104 : 00000;
15105 : 00000;
15106 : 00000;
15107 : 00000;
15110 : 00000;
15111 : 00000;
15112 : 00000;
15113 : 00000;
15114 : 00000;
15115 : 00000;
15116 : 00000;
15117 : 00000;
15120 : 00000;
15121 : 00000;
15122 : 00000;
15123 : 00000;
15124 : 00000;
15125 : 00000;
15126 : 00000;
15127 : 00000;
15130 : 00000;
15131 : 00000;
15132 : 00000;
15133 : 00000;
15134 : 00000;
15135 : 00000;
15136 : 00000;
15137 : 00000;
15140 : 00000;
15141 : 00000;
15142 : 00000;
15143 : 00000;
15144 : 00000;
15145 : 00000;
15146 : 00000;
15147 : 00000;
15150 : 00000;
15151 : 00000;
15152 : 00000;
15153 : 00000;
15154 : 00000;
15155 : 00000;
15156 : 00000;
15157 : 00000;
15160 : 00000;
15161 : 00000;
15162 : 00000;
15163 : 00000;
15164 : 00000;
15165 : 00000;
15166 : 00000;
15167 : 00000;
15170 : 00000;
15171 : 00000;
15172 : 00000;
15173 : 00000;
15174 : 00000;
15175 : 00000;
15176 : 00000;
15177 : 00000;
15200 : 00000;
15201 : 00000;
15202 : 00000;
15203 : 00000;
15204 : 00000;
15205 : 00000;
15206 : 00000;
15207 : 00000;
15210 : 00000;
15211 : 00000;
15212 : 00000;
15213 : 00000;
15214 : 00000;
15215 : 00000;
15216 : 00000;
15217 : 00000;
15220 : 00000;
15221 : 00000;
15222 : 00000;
15223 : 00000;
15224 : 00000;
15225 : 00000;
15226 : 00000;
15227 : 00000;
15230 : 00000;
15231 : 00000;
15232 : 00000;
15233 : 00000;
15234 : 00000;
15235 : 00000;
15236 : 00000;
15237 : 00000;
15240 : 00000;
15241 : 00000;
15242 : 00000;
15243 : 00000;
15244 : 00000;
15245 : 00000;
15246 : 00000;
15247 : 00000;
15250 : 00000;
15251 : 00000;
15252 : 00000;
15253 : 00000;
15254 : 00000;
15255 : 00000;
15256 : 00000;
15257 : 00000;
15260 : 00000;
15261 : 00000;
15262 : 00000;
15263 : 00000;
15264 : 00000;
15265 : 00000;
15266 : 00000;
15267 : 00000;
15270 : 00000;
15271 : 00000;
15272 : 00000;
15273 : 00000;
15274 : 00000;
15275 : 00000;
15276 : 00000;
15277 : 00000;
15300 : 00000;
15301 : 00000;
15302 : 00000;
15303 : 00000;
15304 : 00000;
15305 : 00000;
15306 : 00000;
15307 : 00000;
15310 : 00000;
15311 : 00000;
15312 : 00000;
15313 : 00000;
15314 : 00000;
15315 : 00000;
15316 : 00000;
15317 : 00000;
15320 : 00000;
15321 : 00000;
15322 : 00000;
15323 : 00000;
15324 : 00000;
15325 : 00000;
15326 : 00000;
15327 : 00000;
15330 : 00000;
15331 : 00000;
15332 : 00000;
15333 : 00000;
15334 : 00000;
15335 : 00000;
15336 : 00000;
15337 : 00000;
15340 : 00000;
15341 : 00000;
15342 : 00000;
15343 : 00000;
15344 : 00000;
15345 : 00000;
15346 : 00000;
15347 : 00000;
15350 : 00000;
15351 : 00000;
15352 : 00000;
15353 : 00000;
15354 : 00000;
15355 : 00000;
15356 : 00000;
15357 : 00000;
15360 : 00000;
15361 : 00000;
15362 : 00000;
15363 : 00000;
15364 : 00000;
15365 : 00000;
15366 : 00000;
15367 : 00000;
15370 : 00000;
15371 : 00000;
15372 : 00000;
15373 : 00000;
15374 : 00000;
15375 : 00000;
15376 : 00000;
15377 : 00000;
15400 : 00000;
15401 : 00000;
15402 : 00000;
15403 : 00000;
15404 : 00000;
15405 : 00000;
15406 : 00000;
15407 : 00000;
15410 : 00000;
15411 : 00000;
15412 : 00000;
15413 : 00000;
15414 : 00000;
15415 : 00000;
15416 : 00000;
15417 : 00000;
15420 : 00000;
15421 : 00000;
15422 : 00000;
15423 : 00000;
15424 : 00000;
15425 : 00000;
15426 : 00000;
15427 : 00000;
15430 : 00000;
15431 : 00000;
15432 : 00000;
15433 : 00000;
15434 : 00000;
15435 : 00000;
15436 : 00000;
15437 : 00000;
15440 : 00000;
15441 : 00000;
15442 : 00000;
15443 : 00000;
15444 : 00000;
15445 : 00000;
15446 : 00000;
15447 : 00000;
15450 : 00000;
15451 : 00000;
15452 : 00000;
15453 : 00000;
15454 : 00000;
15455 : 00000;
15456 : 00000;
15457 : 00000;
15460 : 00000;
15461 : 00000;
15462 : 00000;
15463 : 00000;
15464 : 00000;
15465 : 00000;
15466 : 00000;
15467 : 00000;
15470 : 00000;
15471 : 00000;
15472 : 00000;
15473 : 00000;
15474 : 00000;
15475 : 00000;
15476 : 00000;
15477 : 00000;
15500 : 00000;
15501 : 00000;
15502 : 00000;
15503 : 00000;
15504 : 00000;
15505 : 00000;
15506 : 00000;
15507 : 00000;
15510 : 00000;
15511 : 00000;
15512 : 00000;
15513 : 00000;
15514 : 00000;
15515 : 00000;
15516 : 00000;
15517 : 00000;
15520 : 00000;
15521 : 00000;
15522 : 00000;
15523 : 00000;
15524 : 00000;
15525 : 00000;
15526 : 00000;
15527 : 00000;
15530 : 00000;
15531 : 00000;
15532 : 00000;
15533 : 00000;
15534 : 00000;
15535 : 00000;
15536 : 00000;
15537 : 00000;
15540 : 00000;
15541 : 00000;
15542 : 00000;
15543 : 00000;
15544 : 00000;
15545 : 00000;
15546 : 00000;
15547 : 00000;
15550 : 00000;
15551 : 00000;
15552 : 00000;
15553 : 00000;
15554 : 00000;
15555 : 00000;
15556 : 00000;
15557 : 00000;
15560 : 00000;
15561 : 00000;
15562 : 00000;
15563 : 00000;
15564 : 00000;
15565 : 00000;
15566 : 00000;
15567 : 00000;
15570 : 00000;
15571 : 00000;
15572 : 00000;
15573 : 00000;
15574 : 00000;
15575 : 00000;
15576 : 00000;
15577 : 00000;
15600 : 00000;
15601 : 00000;
15602 : 00000;
15603 : 00000;
15604 : 00000;
15605 : 00000;
15606 : 00000;
15607 : 00000;
15610 : 00000;
15611 : 00000;
15612 : 00000;
15613 : 00000;
15614 : 00000;
15615 : 00000;
15616 : 00000;
15617 : 00000;
15620 : 00000;
15621 : 00000;
15622 : 00000;
15623 : 00000;
15624 : 00000;
15625 : 00000;
15626 : 00000;
15627 : 00000;
15630 : 00000;
15631 : 00000;
15632 : 00000;
15633 : 00000;
15634 : 00000;
15635 : 00000;
15636 : 00000;
15637 : 00000;
15640 : 00000;
15641 : 00000;
15642 : 00000;
15643 : 00000;
15644 : 00000;
15645 : 00000;
15646 : 00000;
15647 : 00000;
15650 : 00000;
15651 : 00000;
15652 : 00000;
15653 : 00000;
15654 : 00000;
15655 : 00000;
15656 : 00000;
15657 : 00000;
15660 : 00000;
15661 : 00000;
15662 : 00000;
15663 : 00000;
15664 : 00000;
15665 : 00000;
15666 : 00000;
15667 : 00000;
15670 : 00000;
15671 : 00000;
15672 : 00000;
15673 : 00000;
15674 : 00000;
15675 : 00000;
15676 : 00000;
15677 : 00000;
15700 : 00000;
15701 : 00000;
15702 : 00000;
15703 : 00000;
15704 : 00000;
15705 : 00000;
15706 : 00000;
15707 : 00000;
15710 : 00000;
15711 : 00000;
15712 : 00000;
15713 : 00000;
15714 : 00000;
15715 : 00000;
15716 : 00000;
15717 : 00000;
15720 : 00000;
15721 : 00000;
15722 : 00000;
15723 : 00000;
15724 : 00000;
15725 : 00000;
15726 : 00000;
15727 : 00000;
15730 : 00000;
15731 : 00000;
15732 : 00000;
15733 : 00000;
15734 : 00000;
15735 : 00000;
15736 : 00000;
15737 : 00000;
15740 : 00000;
15741 : 00000;
15742 : 00000;
15743 : 00000;
15744 : 00000;
15745 : 00000;
15746 : 00000;
15747 : 00000;
15750 : 00000;
15751 : 00000;
15752 : 00000;
15753 : 00000;
15754 : 00000;
15755 : 00000;
15756 : 00000;
15757 : 00000;
15760 : 00000;
15761 : 00000;
15762 : 00000;
15763 : 00000;
15764 : 00000;
15765 : 00000;
15766 : 00000;
15767 : 00000;
15770 : 00000;
15771 : 00000;
15772 : 00000;
15773 : 00000;
15774 : 00000;
15775 : 00000;
15776 : 00000;
15777 : 00000;
16000 : 00000;
16001 : 00000;
16002 : 00000;
16003 : 00000;
16004 : 00000;
16005 : 00000;
16006 : 00000;
16007 : 00000;
16010 : 00000;
16011 : 00000;
16012 : 00000;
16013 : 00000;
16014 : 00000;
16015 : 00000;
16016 : 00000;
16017 : 00000;
16020 : 00000;
16021 : 00000;
16022 : 00000;
16023 : 00000;
16024 : 00000;
16025 : 00000;
16026 : 00000;
16027 : 00000;
16030 : 00000;
16031 : 00000;
16032 : 00000;
16033 : 00000;
16034 : 00000;
16035 : 00000;
16036 : 00000;
16037 : 00000;
16040 : 00000;
16041 : 00000;
16042 : 00000;
16043 : 00000;
16044 : 00000;
16045 : 00000;
16046 : 00000;
16047 : 00000;
16050 : 00000;
16051 : 00000;
16052 : 00000;
16053 : 00000;
16054 : 00000;
16055 : 00000;
16056 : 00000;
16057 : 00000;
16060 : 00000;
16061 : 00000;
16062 : 00000;
16063 : 00000;
16064 : 00000;
16065 : 00000;
16066 : 00000;
16067 : 00000;
16070 : 00000;
16071 : 00000;
16072 : 00000;
16073 : 00000;
16074 : 00000;
16075 : 00000;
16076 : 00000;
16077 : 00000;
16100 : 00000;
16101 : 00000;
16102 : 00000;
16103 : 00000;
16104 : 00000;
16105 : 00000;
16106 : 00000;
16107 : 00000;
16110 : 00000;
16111 : 00000;
16112 : 00000;
16113 : 00000;
16114 : 00000;
16115 : 00000;
16116 : 00000;
16117 : 00000;
16120 : 00000;
16121 : 00000;
16122 : 00000;
16123 : 00000;
16124 : 00000;
16125 : 00000;
16126 : 00000;
16127 : 00000;
16130 : 00000;
16131 : 00000;
16132 : 00000;
16133 : 00000;
16134 : 00000;
16135 : 00000;
16136 : 00000;
16137 : 00000;
16140 : 00000;
16141 : 00000;
16142 : 00000;
16143 : 00000;
16144 : 00000;
16145 : 00000;
16146 : 00000;
16147 : 00000;
16150 : 00000;
16151 : 00000;
16152 : 00000;
16153 : 00000;
16154 : 00000;
16155 : 00000;
16156 : 00000;
16157 : 00000;
16160 : 00000;
16161 : 00000;
16162 : 00000;
16163 : 00000;
16164 : 00000;
16165 : 00000;
16166 : 00000;
16167 : 00000;
16170 : 00000;
16171 : 00000;
16172 : 00000;
16173 : 00000;
16174 : 00000;
16175 : 00000;
16176 : 00000;
16177 : 00000;
16200 : 00000;
16201 : 00000;
16202 : 00000;
16203 : 00000;
16204 : 00000;
16205 : 00000;
16206 : 00000;
16207 : 00000;
16210 : 00000;
16211 : 00000;
16212 : 00000;
16213 : 00000;
16214 : 00000;
16215 : 00000;
16216 : 00000;
16217 : 00000;
16220 : 00000;
16221 : 00000;
16222 : 00000;
16223 : 00000;
16224 : 00000;
16225 : 00000;
16226 : 00000;
16227 : 00000;
16230 : 00000;
16231 : 00000;
16232 : 00000;
16233 : 00000;
16234 : 00000;
16235 : 00000;
16236 : 00000;
16237 : 00000;
16240 : 00000;
16241 : 00000;
16242 : 00000;
16243 : 00000;
16244 : 00000;
16245 : 00000;
16246 : 00000;
16247 : 00000;
16250 : 00000;
16251 : 00000;
16252 : 00000;
16253 : 00000;
16254 : 00000;
16255 : 00000;
16256 : 00000;
16257 : 00000;
16260 : 00000;
16261 : 00000;
16262 : 00000;
16263 : 00000;
16264 : 00000;
16265 : 00000;
16266 : 00000;
16267 : 00000;
16270 : 00000;
16271 : 00000;
16272 : 00000;
16273 : 00000;
16274 : 00000;
16275 : 00000;
16276 : 00000;
16277 : 00000;
16300 : 00000;
16301 : 00000;
16302 : 00000;
16303 : 00000;
16304 : 00000;
16305 : 00000;
16306 : 00000;
16307 : 00000;
16310 : 00000;
16311 : 00000;
16312 : 00000;
16313 : 00000;
16314 : 00000;
16315 : 00000;
16316 : 00000;
16317 : 00000;
16320 : 00000;
16321 : 00000;
16322 : 00000;
16323 : 00000;
16324 : 00000;
16325 : 00000;
16326 : 00000;
16327 : 00000;
16330 : 00000;
16331 : 00000;
16332 : 00000;
16333 : 00000;
16334 : 00000;
16335 : 00000;
16336 : 00000;
16337 : 00000;
16340 : 00000;
16341 : 00000;
16342 : 00000;
16343 : 00000;
16344 : 00000;
16345 : 00000;
16346 : 00000;
16347 : 00000;
16350 : 00000;
16351 : 00000;
16352 : 00000;
16353 : 00000;
16354 : 00000;
16355 : 00000;
16356 : 00000;
16357 : 00000;
16360 : 00000;
16361 : 00000;
16362 : 00000;
16363 : 00000;
16364 : 00000;
16365 : 00000;
16366 : 00000;
16367 : 00000;
16370 : 00000;
16371 : 00000;
16372 : 00000;
16373 : 00000;
16374 : 00000;
16375 : 00000;
16376 : 00000;
16377 : 00000;
16400 : 00000;
16401 : 00000;
16402 : 00000;
16403 : 00000;
16404 : 00000;
16405 : 00000;
16406 : 00000;
16407 : 00000;
16410 : 00000;
16411 : 00000;
16412 : 00000;
16413 : 00000;
16414 : 00000;
16415 : 00000;
16416 : 00000;
16417 : 00000;
16420 : 00000;
16421 : 00000;
16422 : 00000;
16423 : 00000;
16424 : 00000;
16425 : 00000;
16426 : 00000;
16427 : 00000;
16430 : 00000;
16431 : 00000;
16432 : 00000;
16433 : 00000;
16434 : 00000;
16435 : 00000;
16436 : 00000;
16437 : 00000;
16440 : 00000;
16441 : 00000;
16442 : 00000;
16443 : 00000;
16444 : 00000;
16445 : 00000;
16446 : 00000;
16447 : 00000;
16450 : 00000;
16451 : 00000;
16452 : 00000;
16453 : 00000;
16454 : 00000;
16455 : 00000;
16456 : 00000;
16457 : 00000;
16460 : 00000;
16461 : 00000;
16462 : 00000;
16463 : 00000;
16464 : 00000;
16465 : 00000;
16466 : 00000;
16467 : 00000;
16470 : 00000;
16471 : 00000;
16472 : 00000;
16473 : 00000;
16474 : 00000;
16475 : 00000;
16476 : 00000;
16477 : 00000;
16500 : 00000;
16501 : 00000;
16502 : 00000;
16503 : 00000;
16504 : 00000;
16505 : 00000;
16506 : 00000;
16507 : 00000;
16510 : 00000;
16511 : 00000;
16512 : 00000;
16513 : 00000;
16514 : 00000;
16515 : 00000;
16516 : 00000;
16517 : 00000;
16520 : 00000;
16521 : 00000;
16522 : 00000;
16523 : 00000;
16524 : 00000;
16525 : 00000;
16526 : 00000;
16527 : 00000;
16530 : 00000;
16531 : 00000;
16532 : 00000;
16533 : 00000;
16534 : 00000;
16535 : 00000;
16536 : 00000;
16537 : 00000;
16540 : 00000;
16541 : 00000;
16542 : 00000;
16543 : 00000;
16544 : 00000;
16545 : 00000;
16546 : 00000;
16547 : 00000;
16550 : 00000;
16551 : 00000;
16552 : 00000;
16553 : 00000;
16554 : 00000;
16555 : 00000;
16556 : 00000;
16557 : 00000;
16560 : 00000;
16561 : 00000;
16562 : 00000;
16563 : 00000;
16564 : 00000;
16565 : 00000;
16566 : 00000;
16567 : 00000;
16570 : 00000;
16571 : 00000;
16572 : 00000;
16573 : 00000;
16574 : 00000;
16575 : 00000;
16576 : 00000;
16577 : 00000;
16600 : 00000;
16601 : 00000;
16602 : 00000;
16603 : 00000;
16604 : 00000;
16605 : 00000;
16606 : 00000;
16607 : 00000;
16610 : 00000;
16611 : 00000;
16612 : 00000;
16613 : 00000;
16614 : 00000;
16615 : 00000;
16616 : 00000;
16617 : 00000;
16620 : 00000;
16621 : 00000;
16622 : 00000;
16623 : 00000;
16624 : 00000;
16625 : 00000;
16626 : 00000;
16627 : 00000;
16630 : 00000;
16631 : 00000;
16632 : 00000;
16633 : 00000;
16634 : 00000;
16635 : 00000;
16636 : 00000;
16637 : 00000;
16640 : 00000;
16641 : 00000;
16642 : 00000;
16643 : 00000;
16644 : 00000;
16645 : 00000;
16646 : 00000;
16647 : 00000;
16650 : 00000;
16651 : 00000;
16652 : 00000;
16653 : 00000;
16654 : 00000;
16655 : 00000;
16656 : 00000;
16657 : 00000;
16660 : 00000;
16661 : 00000;
16662 : 00000;
16663 : 00000;
16664 : 00000;
16665 : 00000;
16666 : 00000;
16667 : 00000;
16670 : 00000;
16671 : 00000;
16672 : 00000;
16673 : 00000;
16674 : 00000;
16675 : 00000;
16676 : 00000;
16677 : 00000;
16700 : 00000;
16701 : 00000;
16702 : 00000;
16703 : 00000;
16704 : 00000;
16705 : 00000;
16706 : 00000;
16707 : 00000;
16710 : 00000;
16711 : 00000;
16712 : 00000;
16713 : 00000;
16714 : 00000;
16715 : 00000;
16716 : 00000;
16717 : 00000;
16720 : 00000;
16721 : 00000;
16722 : 00000;
16723 : 00000;
16724 : 00000;
16725 : 00000;
16726 : 00000;
16727 : 00000;
16730 : 00000;
16731 : 00000;
16732 : 00000;
16733 : 00000;
16734 : 00000;
16735 : 00000;
16736 : 00000;
16737 : 00000;
16740 : 00000;
16741 : 00000;
16742 : 00000;
16743 : 00000;
16744 : 00000;
16745 : 00000;
16746 : 00000;
16747 : 00000;
16750 : 00000;
16751 : 00000;
16752 : 00000;
16753 : 00000;
16754 : 00000;
16755 : 00000;
16756 : 00000;
16757 : 00000;
16760 : 00000;
16761 : 00000;
16762 : 00000;
16763 : 00000;
16764 : 00000;
16765 : 00000;
16766 : 00000;
16767 : 00000;
16770 : 00000;
16771 : 00000;
16772 : 00000;
16773 : 00000;
16774 : 00000;
16775 : 00000;
16776 : 00000;
16777 : 00000;
17000 : 00000;
17001 : 00000;
17002 : 00000;
17003 : 00000;
17004 : 00000;
17005 : 00000;
17006 : 00000;
17007 : 00000;
17010 : 00000;
17011 : 00000;
17012 : 00000;
17013 : 00000;
17014 : 00000;
17015 : 00000;
17016 : 00000;
17017 : 00000;
17020 : 00000;
17021 : 00000;
17022 : 00000;
17023 : 00000;
17024 : 00000;
17025 : 00000;
17026 : 00000;
17027 : 00000;
17030 : 00000;
17031 : 00000;
17032 : 00000;
17033 : 00000;
17034 : 00000;
17035 : 00000;
17036 : 00000;
17037 : 00000;
17040 : 00000;
17041 : 00000;
17042 : 00000;
17043 : 00000;
17044 : 00000;
17045 : 00000;
17046 : 00000;
17047 : 00000;
17050 : 00000;
17051 : 00000;
17052 : 00000;
17053 : 00000;
17054 : 00000;
17055 : 00000;
17056 : 00000;
17057 : 00000;
17060 : 00000;
17061 : 00000;
17062 : 00000;
17063 : 00000;
17064 : 00000;
17065 : 00000;
17066 : 00000;
17067 : 00000;
17070 : 00000;
17071 : 00000;
17072 : 00000;
17073 : 00000;
17074 : 00000;
17075 : 00000;
17076 : 00000;
17077 : 00000;
17100 : 00000;
17101 : 00000;
17102 : 00000;
17103 : 00000;
17104 : 00000;
17105 : 00000;
17106 : 00000;
17107 : 00000;
17110 : 00000;
17111 : 00000;
17112 : 00000;
17113 : 00000;
17114 : 00000;
17115 : 00000;
17116 : 00000;
17117 : 00000;
17120 : 00000;
17121 : 00000;
17122 : 00000;
17123 : 00000;
17124 : 00000;
17125 : 00000;
17126 : 00000;
17127 : 00000;
17130 : 00000;
17131 : 00000;
17132 : 00000;
17133 : 00000;
17134 : 00000;
17135 : 00000;
17136 : 00000;
17137 : 00000;
17140 : 00000;
17141 : 00000;
17142 : 00000;
17143 : 00000;
17144 : 00000;
17145 : 00000;
17146 : 00000;
17147 : 00000;
17150 : 00000;
17151 : 00000;
17152 : 00000;
17153 : 00000;
17154 : 00000;
17155 : 00000;
17156 : 00000;
17157 : 00000;
17160 : 00000;
17161 : 00000;
17162 : 00000;
17163 : 00000;
17164 : 00000;
17165 : 00000;
17166 : 00000;
17167 : 00000;
17170 : 00000;
17171 : 00000;
17172 : 00000;
17173 : 00000;
17174 : 00000;
17175 : 00000;
17176 : 00000;
17177 : 00000;
17200 : 00000;
17201 : 00000;
17202 : 00000;
17203 : 00000;
17204 : 00000;
17205 : 00000;
17206 : 00000;
17207 : 00000;
17210 : 00000;
17211 : 00000;
17212 : 00000;
17213 : 00000;
17214 : 00000;
17215 : 00000;
17216 : 00000;
17217 : 00000;
17220 : 00000;
17221 : 00000;
17222 : 00000;
17223 : 00000;
17224 : 00000;
17225 : 00000;
17226 : 00000;
17227 : 00000;
17230 : 00000;
17231 : 00000;
17232 : 00000;
17233 : 00000;
17234 : 00000;
17235 : 00000;
17236 : 00000;
17237 : 00000;
17240 : 00000;
17241 : 00000;
17242 : 00000;
17243 : 00000;
17244 : 00000;
17245 : 00000;
17246 : 00000;
17247 : 00000;
17250 : 00000;
17251 : 00000;
17252 : 00000;
17253 : 00000;
17254 : 00000;
17255 : 00000;
17256 : 00000;
17257 : 00000;
17260 : 00000;
17261 : 00000;
17262 : 00000;
17263 : 00000;
17264 : 00000;
17265 : 00000;
17266 : 00000;
17267 : 00000;
17270 : 00000;
17271 : 00000;
17272 : 00000;
17273 : 00000;
17274 : 00000;
17275 : 00000;
17276 : 00000;
17277 : 00000;
17300 : 00000;
17301 : 00000;
17302 : 00000;
17303 : 00000;
17304 : 00000;
17305 : 00000;
17306 : 00000;
17307 : 00000;
17310 : 00000;
17311 : 00000;
17312 : 00000;
17313 : 00000;
17314 : 00000;
17315 : 00000;
17316 : 00000;
17317 : 00000;
17320 : 00000;
17321 : 00000;
17322 : 00000;
17323 : 00000;
17324 : 00000;
17325 : 00000;
17326 : 00000;
17327 : 00000;
17330 : 00000;
17331 : 00000;
17332 : 00000;
17333 : 00000;
17334 : 00000;
17335 : 00000;
17336 : 00000;
17337 : 00000;
17340 : 00000;
17341 : 00000;
17342 : 00000;
17343 : 00000;
17344 : 00000;
17345 : 00000;
17346 : 00000;
17347 : 00000;
17350 : 00000;
17351 : 00000;
17352 : 00000;
17353 : 00000;
17354 : 00000;
17355 : 00000;
17356 : 00000;
17357 : 00000;
17360 : 00000;
17361 : 00000;
17362 : 00000;
17363 : 00000;
17364 : 00000;
17365 : 00000;
17366 : 00000;
17367 : 00000;
17370 : 00000;
17371 : 00000;
17372 : 00000;
17373 : 00000;
17374 : 00000;
17375 : 00000;
17376 : 00000;
17377 : 00000;
17400 : 00000;
17401 : 00000;
17402 : 00000;
17403 : 00000;
17404 : 00000;
17405 : 00000;
17406 : 00000;
17407 : 00000;
17410 : 00000;
17411 : 00000;
17412 : 00000;
17413 : 00000;
17414 : 00000;
17415 : 00000;
17416 : 00000;
17417 : 00000;
17420 : 00000;
17421 : 00000;
17422 : 00000;
17423 : 00000;
17424 : 00000;
17425 : 00000;
17426 : 00000;
17427 : 00000;
17430 : 00000;
17431 : 00000;
17432 : 00000;
17433 : 00000;
17434 : 00000;
17435 : 00000;
17436 : 00000;
17437 : 00000;
17440 : 00000;
17441 : 00000;
17442 : 00000;
17443 : 00000;
17444 : 00000;
17445 : 00000;
17446 : 00000;
17447 : 00000;
17450 : 00000;
17451 : 00000;
17452 : 00000;
17453 : 00000;
17454 : 00000;
17455 : 00000;
17456 : 00000;
17457 : 00000;
17460 : 00000;
17461 : 00000;
17462 : 00000;
17463 : 00000;
17464 : 00000;
17465 : 00000;
17466 : 00000;
17467 : 00000;
17470 : 00000;
17471 : 00000;
17472 : 00000;
17473 : 00000;
17474 : 00000;
17475 : 00000;
17476 : 00000;
17477 : 00000;
17500 : 00000;
17501 : 00000;
17502 : 00000;
17503 : 00000;
17504 : 00000;
17505 : 00000;
17506 : 00000;
17507 : 00000;
17510 : 00000;
17511 : 00000;
17512 : 00000;
17513 : 00000;
17514 : 00000;
17515 : 00000;
17516 : 00000;
17517 : 00000;
17520 : 00000;
17521 : 00000;
17522 : 00000;
17523 : 00000;
17524 : 00000;
17525 : 00000;
17526 : 00000;
17527 : 00000;
17530 : 00000;
17531 : 00000;
17532 : 00000;
17533 : 00000;
17534 : 00000;
17535 : 00000;
17536 : 00000;
17537 : 00000;
17540 : 00000;
17541 : 00000;
17542 : 00000;
17543 : 00000;
17544 : 00000;
17545 : 00000;
17546 : 00000;
17547 : 00000;
17550 : 00000;
17551 : 00000;
17552 : 00000;
17553 : 00000;
17554 : 00000;
17555 : 00000;
17556 : 00000;
17557 : 00000;
17560 : 00000;
17561 : 00000;
17562 : 00000;
17563 : 00000;
17564 : 00000;
17565 : 00000;
17566 : 00000;
17567 : 00000;
17570 : 00000;
17571 : 00000;
17572 : 00000;
17573 : 00000;
17574 : 00000;
17575 : 00000;
17576 : 00000;
17577 : 00000;
17600 : 00000;
17601 : 00000;
17602 : 00000;
17603 : 00000;
17604 : 00000;
17605 : 00000;
17606 : 00000;
17607 : 00000;
17610 : 00000;
17611 : 00000;
17612 : 00000;
17613 : 00000;
17614 : 00000;
17615 : 00000;
17616 : 00000;
17617 : 00000;
17620 : 00000;
17621 : 00000;
17622 : 00000;
17623 : 00000;
17624 : 00000;
17625 : 00000;
17626 : 00000;
17627 : 00000;
17630 : 00000;
17631 : 00000;
17632 : 00000;
17633 : 00000;
17634 : 00000;
17635 : 00000;
17636 : 00000;
17637 : 00000;
17640 : 00000;
17641 : 00000;
17642 : 00000;
17643 : 00000;
17644 : 00000;
17645 : 00000;
17646 : 00000;
17647 : 00000;
17650 : 00000;
17651 : 00000;
17652 : 00000;
17653 : 00000;
17654 : 00000;
17655 : 00000;
17656 : 00000;
17657 : 00000;
17660 : 00000;
17661 : 00000;
17662 : 00000;
17663 : 00000;
17664 : 00000;
17665 : 00000;
17666 : 00000;
17667 : 00000;
17670 : 00000;
17671 : 00000;
17672 : 00000;
17673 : 00000;
17674 : 00000;
17675 : 00000;
17676 : 00000;
17677 : 00000;
17700 : 00000;
17701 : 00000;
17702 : 00000;
17703 : 00000;
17704 : 00000;
17705 : 00000;
17706 : 00000;
17707 : 00000;
17710 : 00000;
17711 : 00000;
17712 : 00000;
17713 : 00000;
17714 : 00000;
17715 : 00000;
17716 : 00000;
17717 : 00000;
17720 : 00000;
17721 : 00000;
17722 : 00000;
17723 : 00000;
17724 : 00000;
17725 : 00000;
17726 : 00000;
17727 : 00000;
17730 : 00000;
17731 : 00000;
17732 : 00000;
17733 : 00000;
17734 : 00000;
17735 : 00000;
17736 : 00000;
17737 : 00000;
17740 : 00000;
17741 : 00000;
17742 : 00000;
17743 : 00000;
17744 : 00000;
17745 : 00000;
17746 : 00000;
17747 : 00000;
17750 : 00000;
17751 : 00000;
17752 : 00000;
17753 : 00000;
17754 : 00000;
17755 : 00000;
17756 : 00000;
17757 : 00000;
17760 : 00000;
17761 : 00000;
17762 : 00000;
17763 : 00000;
17764 : 00000;
17765 : 00000;
17766 : 00000;
17767 : 00000;
17770 : 00000;
17771 : 00000;
17772 : 00000;
17773 : 00000;
17774 : 00000;
17775 : 00000;
17776 : 00000;
17777 : 00000;
20000 : 00000;
20001 : 00000;
20002 : 00000;
20003 : 00000;
20004 : 00000;
20005 : 00000;
20006 : 00000;
20007 : 00000;
20010 : 00000;
20011 : 00000;
20012 : 00000;
20013 : 00000;
20014 : 00000;
20015 : 00000;
20016 : 00000;
20017 : 00000;
20020 : 00000;
20021 : 00000;
20022 : 00000;
20023 : 00000;
20024 : 00000;
20025 : 00000;
20026 : 00000;
20027 : 00000;
20030 : 00000;
20031 : 00000;
20032 : 00000;
20033 : 00000;
20034 : 00000;
20035 : 00000;
20036 : 00000;
20037 : 00000;
20040 : 00000;
20041 : 00000;
20042 : 00000;
20043 : 00000;
20044 : 00000;
20045 : 00000;
20046 : 00000;
20047 : 00000;
20050 : 00000;
20051 : 00000;
20052 : 00000;
20053 : 00000;
20054 : 00000;
20055 : 00000;
20056 : 00000;
20057 : 00000;
20060 : 00000;
20061 : 00000;
20062 : 00000;
20063 : 00000;
20064 : 00000;
20065 : 00000;
20066 : 00000;
20067 : 00000;
20070 : 00000;
20071 : 00000;
20072 : 00000;
20073 : 00000;
20074 : 00000;
20075 : 00000;
20076 : 00000;
20077 : 00000;
20100 : 00000;
20101 : 00000;
20102 : 00000;
20103 : 00000;
20104 : 00000;
20105 : 00000;
20106 : 00000;
20107 : 00000;
20110 : 00000;
20111 : 00000;
20112 : 00000;
20113 : 00000;
20114 : 00000;
20115 : 00000;
20116 : 00000;
20117 : 00000;
20120 : 00000;
20121 : 00000;
20122 : 00000;
20123 : 00000;
20124 : 00000;
20125 : 00000;
20126 : 00000;
20127 : 00000;
20130 : 00000;
20131 : 00000;
20132 : 00000;
20133 : 00000;
20134 : 00000;
20135 : 00000;
20136 : 00000;
20137 : 00000;
20140 : 00000;
20141 : 00000;
20142 : 00000;
20143 : 00000;
20144 : 00000;
20145 : 00000;
20146 : 00000;
20147 : 00000;
20150 : 00000;
20151 : 00000;
20152 : 00000;
20153 : 00000;
20154 : 00000;
20155 : 00000;
20156 : 00000;
20157 : 00000;
20160 : 00000;
20161 : 00000;
20162 : 00000;
20163 : 00000;
20164 : 00000;
20165 : 00000;
20166 : 00000;
20167 : 00000;
20170 : 00000;
20171 : 00000;
20172 : 00000;
20173 : 00000;
20174 : 00000;
20175 : 00000;
20176 : 00000;
20177 : 00000;
20200 : 00000;
20201 : 00000;
20202 : 00000;
20203 : 00000;
20204 : 00000;
20205 : 00000;
20206 : 00000;
20207 : 00000;
20210 : 00000;
20211 : 00000;
20212 : 00000;
20213 : 00000;
20214 : 00000;
20215 : 00000;
20216 : 00000;
20217 : 00000;
20220 : 00000;
20221 : 00000;
20222 : 00000;
20223 : 00000;
20224 : 00000;
20225 : 00000;
20226 : 00000;
20227 : 00000;
20230 : 00000;
20231 : 00000;
20232 : 00000;
20233 : 00000;
20234 : 00000;
20235 : 00000;
20236 : 00000;
20237 : 00000;
20240 : 00000;
20241 : 00000;
20242 : 00000;
20243 : 00000;
20244 : 00000;
20245 : 00000;
20246 : 00000;
20247 : 00000;
20250 : 00000;
20251 : 00000;
20252 : 00000;
20253 : 00000;
20254 : 00000;
20255 : 00000;
20256 : 00000;
20257 : 00000;
20260 : 00000;
20261 : 00000;
20262 : 00000;
20263 : 00000;
20264 : 00000;
20265 : 00000;
20266 : 00000;
20267 : 00000;
20270 : 00000;
20271 : 00000;
20272 : 00000;
20273 : 00000;
20274 : 00000;
20275 : 00000;
20276 : 00000;
20277 : 00000;
20300 : 00000;
20301 : 00000;
20302 : 00000;
20303 : 00000;
20304 : 00000;
20305 : 00000;
20306 : 00000;
20307 : 00000;
20310 : 00000;
20311 : 00000;
20312 : 00000;
20313 : 00000;
20314 : 00000;
20315 : 00000;
20316 : 00000;
20317 : 00000;
20320 : 00000;
20321 : 00000;
20322 : 00000;
20323 : 00000;
20324 : 00000;
20325 : 00000;
20326 : 00000;
20327 : 00000;
20330 : 00000;
20331 : 00000;
20332 : 00000;
20333 : 00000;
20334 : 00000;
20335 : 00000;
20336 : 00000;
20337 : 00000;
20340 : 00000;
20341 : 00000;
20342 : 00000;
20343 : 00000;
20344 : 00000;
20345 : 00000;
20346 : 00000;
20347 : 00000;
20350 : 00000;
20351 : 00000;
20352 : 00000;
20353 : 00000;
20354 : 00000;
20355 : 00000;
20356 : 00000;
20357 : 00000;
20360 : 00000;
20361 : 00000;
20362 : 00000;
20363 : 00000;
20364 : 00000;
20365 : 00000;
20366 : 00000;
20367 : 00000;
20370 : 00000;
20371 : 00000;
20372 : 00000;
20373 : 00000;
20374 : 00000;
20375 : 00000;
20376 : 00000;
20377 : 00000;
20400 : 00000;
20401 : 00000;
20402 : 00000;
20403 : 00000;
20404 : 00000;
20405 : 00000;
20406 : 00000;
20407 : 00000;
20410 : 00000;
20411 : 00000;
20412 : 00000;
20413 : 00000;
20414 : 00000;
20415 : 00000;
20416 : 00000;
20417 : 00000;
20420 : 00000;
20421 : 00000;
20422 : 00000;
20423 : 00000;
20424 : 00000;
20425 : 00000;
20426 : 00000;
20427 : 00000;
20430 : 00000;
20431 : 00000;
20432 : 00000;
20433 : 00000;
20434 : 00000;
20435 : 00000;
20436 : 00000;
20437 : 00000;
20440 : 00000;
20441 : 00000;
20442 : 00000;
20443 : 00000;
20444 : 00000;
20445 : 00000;
20446 : 00000;
20447 : 00000;
20450 : 00000;
20451 : 00000;
20452 : 00000;
20453 : 00000;
20454 : 00000;
20455 : 00000;
20456 : 00000;
20457 : 00000;
20460 : 00000;
20461 : 00000;
20462 : 00000;
20463 : 00000;
20464 : 00000;
20465 : 00000;
20466 : 00000;
20467 : 00000;
20470 : 00000;
20471 : 00000;
20472 : 00000;
20473 : 00000;
20474 : 00000;
20475 : 00000;
20476 : 00000;
20477 : 00000;
20500 : 00000;
20501 : 00000;
20502 : 00000;
20503 : 00000;
20504 : 00000;
20505 : 00000;
20506 : 00000;
20507 : 00000;
20510 : 00000;
20511 : 00000;
20512 : 00000;
20513 : 00000;
20514 : 00000;
20515 : 00000;
20516 : 00000;
20517 : 00000;
20520 : 00000;
20521 : 00000;
20522 : 00000;
20523 : 00000;
20524 : 00000;
20525 : 00000;
20526 : 00000;
20527 : 00000;
20530 : 00000;
20531 : 00000;
20532 : 00000;
20533 : 00000;
20534 : 00000;
20535 : 00000;
20536 : 00000;
20537 : 00000;
20540 : 00000;
20541 : 00000;
20542 : 00000;
20543 : 00000;
20544 : 00000;
20545 : 00000;
20546 : 00000;
20547 : 00000;
20550 : 00000;
20551 : 00000;
20552 : 00000;
20553 : 00000;
20554 : 00000;
20555 : 00000;
20556 : 00000;
20557 : 00000;
20560 : 00000;
20561 : 00000;
20562 : 00000;
20563 : 00000;
20564 : 00000;
20565 : 00000;
20566 : 00000;
20567 : 00000;
20570 : 00000;
20571 : 00000;
20572 : 00000;
20573 : 00000;
20574 : 00000;
20575 : 00000;
20576 : 00000;
20577 : 00000;
20600 : 00000;
20601 : 00000;
20602 : 00000;
20603 : 00000;
20604 : 00000;
20605 : 00000;
20606 : 00000;
20607 : 00000;
20610 : 00000;
20611 : 00000;
20612 : 00000;
20613 : 00000;
20614 : 00000;
20615 : 00000;
20616 : 00000;
20617 : 00000;
20620 : 00000;
20621 : 00000;
20622 : 00000;
20623 : 00000;
20624 : 00000;
20625 : 00000;
20626 : 00000;
20627 : 00000;
20630 : 00000;
20631 : 00000;
20632 : 00000;
20633 : 00000;
20634 : 00000;
20635 : 00000;
20636 : 00000;
20637 : 00000;
20640 : 00000;
20641 : 00000;
20642 : 00000;
20643 : 00000;
20644 : 00000;
20645 : 00000;
20646 : 00000;
20647 : 00000;
20650 : 00000;
20651 : 00000;
20652 : 00000;
20653 : 00000;
20654 : 00000;
20655 : 00000;
20656 : 00000;
20657 : 00000;
20660 : 00000;
20661 : 00000;
20662 : 00000;
20663 : 00000;
20664 : 00000;
20665 : 00000;
20666 : 00000;
20667 : 00000;
20670 : 00000;
20671 : 00000;
20672 : 00000;
20673 : 00000;
20674 : 00000;
20675 : 00000;
20676 : 00000;
20677 : 00000;
20700 : 00000;
20701 : 00000;
20702 : 00000;
20703 : 00000;
20704 : 00000;
20705 : 00000;
20706 : 00000;
20707 : 00000;
20710 : 00000;
20711 : 00000;
20712 : 00000;
20713 : 00000;
20714 : 00000;
20715 : 00000;
20716 : 00000;
20717 : 00000;
20720 : 00000;
20721 : 00000;
20722 : 00000;
20723 : 00000;
20724 : 00000;
20725 : 00000;
20726 : 00000;
20727 : 00000;
20730 : 00000;
20731 : 00000;
20732 : 00000;
20733 : 00000;
20734 : 00000;
20735 : 00000;
20736 : 00000;
20737 : 00000;
20740 : 00000;
20741 : 00000;
20742 : 00000;
20743 : 00000;
20744 : 00000;
20745 : 00000;
20746 : 00000;
20747 : 00000;
20750 : 00000;
20751 : 00000;
20752 : 00000;
20753 : 00000;
20754 : 00000;
20755 : 00000;
20756 : 00000;
20757 : 00000;
20760 : 00000;
20761 : 00000;
20762 : 00000;
20763 : 00000;
20764 : 00000;
20765 : 00000;
20766 : 00000;
20767 : 00000;
20770 : 00000;
20771 : 00000;
20772 : 00000;
20773 : 00000;
20774 : 00000;
20775 : 00000;
20776 : 00000;
20777 : 00000;
21000 : 00000;
21001 : 00000;
21002 : 00000;
21003 : 00000;
21004 : 00000;
21005 : 00000;
21006 : 00000;
21007 : 00000;
21010 : 00000;
21011 : 00000;
21012 : 00000;
21013 : 00000;
21014 : 00000;
21015 : 00000;
21016 : 00000;
21017 : 00000;
21020 : 00000;
21021 : 00000;
21022 : 00000;
21023 : 00000;
21024 : 00000;
21025 : 00000;
21026 : 00000;
21027 : 00000;
21030 : 00000;
21031 : 00000;
21032 : 00000;
21033 : 00000;
21034 : 00000;
21035 : 00000;
21036 : 00000;
21037 : 00000;
21040 : 00000;
21041 : 00000;
21042 : 00000;
21043 : 00000;
21044 : 00000;
21045 : 00000;
21046 : 00000;
21047 : 00000;
21050 : 00000;
21051 : 00000;
21052 : 00000;
21053 : 00000;
21054 : 00000;
21055 : 00000;
21056 : 00000;
21057 : 00000;
21060 : 00000;
21061 : 00000;
21062 : 00000;
21063 : 00000;
21064 : 00000;
21065 : 00000;
21066 : 00000;
21067 : 00000;
21070 : 00000;
21071 : 00000;
21072 : 00000;
21073 : 00000;
21074 : 00000;
21075 : 00000;
21076 : 00000;
21077 : 00000;
21100 : 00000;
21101 : 00000;
21102 : 00000;
21103 : 00000;
21104 : 00000;
21105 : 00000;
21106 : 00000;
21107 : 00000;
21110 : 00000;
21111 : 00000;
21112 : 00000;
21113 : 00000;
21114 : 00000;
21115 : 00000;
21116 : 00000;
21117 : 00000;
21120 : 00000;
21121 : 00000;
21122 : 00000;
21123 : 00000;
21124 : 00000;
21125 : 00000;
21126 : 00000;
21127 : 00000;
21130 : 00000;
21131 : 00000;
21132 : 00000;
21133 : 00000;
21134 : 00000;
21135 : 00000;
21136 : 00000;
21137 : 00000;
21140 : 00000;
21141 : 00000;
21142 : 00000;
21143 : 00000;
21144 : 00000;
21145 : 00000;
21146 : 00000;
21147 : 00000;
21150 : 00000;
21151 : 00000;
21152 : 00000;
21153 : 00000;
21154 : 00000;
21155 : 00000;
21156 : 00000;
21157 : 00000;
21160 : 00000;
21161 : 00000;
21162 : 00000;
21163 : 00000;
21164 : 00000;
21165 : 00000;
21166 : 00000;
21167 : 00000;
21170 : 00000;
21171 : 00000;
21172 : 00000;
21173 : 00000;
21174 : 00000;
21175 : 00000;
21176 : 00000;
21177 : 00000;
21200 : 00000;
21201 : 00000;
21202 : 00000;
21203 : 00000;
21204 : 00000;
21205 : 00000;
21206 : 00000;
21207 : 00000;
21210 : 00000;
21211 : 00000;
21212 : 00000;
21213 : 00000;
21214 : 00000;
21215 : 00000;
21216 : 00000;
21217 : 00000;
21220 : 00000;
21221 : 00000;
21222 : 00000;
21223 : 00000;
21224 : 00000;
21225 : 00000;
21226 : 00000;
21227 : 00000;
21230 : 00000;
21231 : 00000;
21232 : 00000;
21233 : 00000;
21234 : 00000;
21235 : 00000;
21236 : 00000;
21237 : 00000;
21240 : 00000;
21241 : 00000;
21242 : 00000;
21243 : 00000;
21244 : 00000;
21245 : 00000;
21246 : 00000;
21247 : 00000;
21250 : 00000;
21251 : 00000;
21252 : 00000;
21253 : 00000;
21254 : 00000;
21255 : 00000;
21256 : 00000;
21257 : 00000;
21260 : 00000;
21261 : 00000;
21262 : 00000;
21263 : 00000;
21264 : 00000;
21265 : 00000;
21266 : 00000;
21267 : 00000;
21270 : 00000;
21271 : 00000;
21272 : 00000;
21273 : 00000;
21274 : 00000;
21275 : 00000;
21276 : 00000;
21277 : 00000;
21300 : 00000;
21301 : 00000;
21302 : 00000;
21303 : 00000;
21304 : 00000;
21305 : 00000;
21306 : 00000;
21307 : 00000;
21310 : 00000;
21311 : 00000;
21312 : 00000;
21313 : 00000;
21314 : 00000;
21315 : 00000;
21316 : 00000;
21317 : 00000;
21320 : 00000;
21321 : 00000;
21322 : 00000;
21323 : 00000;
21324 : 00000;
21325 : 00000;
21326 : 00000;
21327 : 00000;
21330 : 00000;
21331 : 00000;
21332 : 00000;
21333 : 00000;
21334 : 00000;
21335 : 00000;
21336 : 00000;
21337 : 00000;
21340 : 00000;
21341 : 00000;
21342 : 00000;
21343 : 00000;
21344 : 00000;
21345 : 00000;
21346 : 00000;
21347 : 00000;
21350 : 00000;
21351 : 00000;
21352 : 00000;
21353 : 00000;
21354 : 00000;
21355 : 00000;
21356 : 00000;
21357 : 00000;
21360 : 00000;
21361 : 00000;
21362 : 00000;
21363 : 00000;
21364 : 00000;
21365 : 00000;
21366 : 00000;
21367 : 00000;
21370 : 00000;
21371 : 00000;
21372 : 00000;
21373 : 00000;
21374 : 00000;
21375 : 00000;
21376 : 00000;
21377 : 00000;
21400 : 00000;
21401 : 00000;
21402 : 00000;
21403 : 00000;
21404 : 00000;
21405 : 00000;
21406 : 00000;
21407 : 00000;
21410 : 00000;
21411 : 00000;
21412 : 00000;
21413 : 00000;
21414 : 00000;
21415 : 00000;
21416 : 00000;
21417 : 00000;
21420 : 00000;
21421 : 00000;
21422 : 00000;
21423 : 00000;
21424 : 00000;
21425 : 00000;
21426 : 00000;
21427 : 00000;
21430 : 00000;
21431 : 00000;
21432 : 00000;
21433 : 00000;
21434 : 00000;
21435 : 00000;
21436 : 00000;
21437 : 00000;
21440 : 00000;
21441 : 00000;
21442 : 00000;
21443 : 00000;
21444 : 00000;
21445 : 00000;
21446 : 00000;
21447 : 00000;
21450 : 00000;
21451 : 00000;
21452 : 00000;
21453 : 00000;
21454 : 00000;
21455 : 00000;
21456 : 00000;
21457 : 00000;
21460 : 00000;
21461 : 00000;
21462 : 00000;
21463 : 00000;
21464 : 00000;
21465 : 00000;
21466 : 00000;
21467 : 00000;
21470 : 00000;
21471 : 00000;
21472 : 00000;
21473 : 00000;
21474 : 00000;
21475 : 00000;
21476 : 00000;
21477 : 00000;
21500 : 00000;
21501 : 00000;
21502 : 00000;
21503 : 00000;
21504 : 00000;
21505 : 00000;
21506 : 00000;
21507 : 00000;
21510 : 00000;
21511 : 00000;
21512 : 00000;
21513 : 00000;
21514 : 00000;
21515 : 00000;
21516 : 00000;
21517 : 00000;
21520 : 00000;
21521 : 00000;
21522 : 00000;
21523 : 00000;
21524 : 00000;
21525 : 00000;
21526 : 00000;
21527 : 00000;
21530 : 00000;
21531 : 00000;
21532 : 00000;
21533 : 00000;
21534 : 00000;
21535 : 00000;
21536 : 00000;
21537 : 00000;
21540 : 00000;
21541 : 00000;
21542 : 00000;
21543 : 00000;
21544 : 00000;
21545 : 00000;
21546 : 00000;
21547 : 00000;
21550 : 00000;
21551 : 00000;
21552 : 00000;
21553 : 00000;
21554 : 00000;
21555 : 00000;
21556 : 00000;
21557 : 00000;
21560 : 00000;
21561 : 00000;
21562 : 00000;
21563 : 00000;
21564 : 00000;
21565 : 00000;
21566 : 00000;
21567 : 00000;
21570 : 00000;
21571 : 00000;
21572 : 00000;
21573 : 00000;
21574 : 00000;
21575 : 00000;
21576 : 00000;
21577 : 00000;
21600 : 00000;
21601 : 00000;
21602 : 00000;
21603 : 00000;
21604 : 00000;
21605 : 00000;
21606 : 00000;
21607 : 00000;
21610 : 00000;
21611 : 00000;
21612 : 00000;
21613 : 00000;
21614 : 00000;
21615 : 00000;
21616 : 00000;
21617 : 00000;
21620 : 00000;
21621 : 00000;
21622 : 00000;
21623 : 00000;
21624 : 00000;
21625 : 00000;
21626 : 00000;
21627 : 00000;
21630 : 00000;
21631 : 00000;
21632 : 00000;
21633 : 00000;
21634 : 00000;
21635 : 00000;
21636 : 00000;
21637 : 00000;
21640 : 00000;
21641 : 00000;
21642 : 00000;
21643 : 00000;
21644 : 00000;
21645 : 00000;
21646 : 00000;
21647 : 00000;
21650 : 00000;
21651 : 00000;
21652 : 00000;
21653 : 00000;
21654 : 00000;
21655 : 00000;
21656 : 00000;
21657 : 00000;
21660 : 00000;
21661 : 00000;
21662 : 00000;
21663 : 00000;
21664 : 00000;
21665 : 00000;
21666 : 00000;
21667 : 00000;
21670 : 00000;
21671 : 00000;
21672 : 00000;
21673 : 00000;
21674 : 00000;
21675 : 00000;
21676 : 00000;
21677 : 00000;
21700 : 00000;
21701 : 00000;
21702 : 00000;
21703 : 00000;
21704 : 00000;
21705 : 00000;
21706 : 00000;
21707 : 00000;
21710 : 00000;
21711 : 00000;
21712 : 00000;
21713 : 00000;
21714 : 00000;
21715 : 00000;
21716 : 00000;
21717 : 00000;
21720 : 00000;
21721 : 00000;
21722 : 00000;
21723 : 00000;
21724 : 00000;
21725 : 00000;
21726 : 00000;
21727 : 00000;
21730 : 00000;
21731 : 00000;
21732 : 00000;
21733 : 00000;
21734 : 00000;
21735 : 00000;
21736 : 00000;
21737 : 00000;
21740 : 00000;
21741 : 00000;
21742 : 00000;
21743 : 00000;
21744 : 00000;
21745 : 00000;
21746 : 00000;
21747 : 00000;
21750 : 00000;
21751 : 00000;
21752 : 00000;
21753 : 00000;
21754 : 00000;
21755 : 00000;
21756 : 00000;
21757 : 00000;
21760 : 00000;
21761 : 00000;
21762 : 00000;
21763 : 00000;
21764 : 00000;
21765 : 00000;
21766 : 00000;
21767 : 00000;
21770 : 00000;
21771 : 00000;
21772 : 00000;
21773 : 00000;
21774 : 00000;
21775 : 00000;
21776 : 00000;
21777 : 00000;
22000 : 00000;
22001 : 00000;
22002 : 00000;
22003 : 00000;
22004 : 00000;
22005 : 00000;
22006 : 00000;
22007 : 00000;
22010 : 00000;
22011 : 00000;
22012 : 00000;
22013 : 00000;
22014 : 00000;
22015 : 00000;
22016 : 00000;
22017 : 00000;
22020 : 00000;
22021 : 00000;
22022 : 00000;
22023 : 00000;
22024 : 00000;
22025 : 00000;
22026 : 00000;
22027 : 00000;
22030 : 00000;
22031 : 00000;
22032 : 00000;
22033 : 00000;
22034 : 00000;
22035 : 00000;
22036 : 00000;
22037 : 00000;
22040 : 00000;
22041 : 00000;
22042 : 00000;
22043 : 00000;
22044 : 00000;
22045 : 00000;
22046 : 00000;
22047 : 00000;
22050 : 00000;
22051 : 00000;
22052 : 00000;
22053 : 00000;
22054 : 00000;
22055 : 00000;
22056 : 00000;
22057 : 00000;
22060 : 00000;
22061 : 00000;
22062 : 00000;
22063 : 00000;
22064 : 00000;
22065 : 00000;
22066 : 00000;
22067 : 00000;
22070 : 00000;
22071 : 00000;
22072 : 00000;
22073 : 00000;
22074 : 00000;
22075 : 00000;
22076 : 00000;
22077 : 00000;
22100 : 00000;
22101 : 00000;
22102 : 00000;
22103 : 00000;
22104 : 00000;
22105 : 00000;
22106 : 00000;
22107 : 00000;
22110 : 00000;
22111 : 00000;
22112 : 00000;
22113 : 00000;
22114 : 00000;
22115 : 00000;
22116 : 00000;
22117 : 00000;
22120 : 00000;
22121 : 00000;
22122 : 00000;
22123 : 00000;
22124 : 00000;
22125 : 00000;
22126 : 00000;
22127 : 00000;
22130 : 00000;
22131 : 00000;
22132 : 00000;
22133 : 00000;
22134 : 00000;
22135 : 00000;
22136 : 00000;
22137 : 00000;
22140 : 00000;
22141 : 00000;
22142 : 00000;
22143 : 00000;
22144 : 00000;
22145 : 00000;
22146 : 00000;
22147 : 00000;
22150 : 00000;
22151 : 00000;
22152 : 00000;
22153 : 00000;
22154 : 00000;
22155 : 00000;
22156 : 00000;
22157 : 00000;
22160 : 00000;
22161 : 00000;
22162 : 00000;
22163 : 00000;
22164 : 00000;
22165 : 00000;
22166 : 00000;
22167 : 00000;
22170 : 00000;
22171 : 00000;
22172 : 00000;
22173 : 00000;
22174 : 00000;
22175 : 00000;
22176 : 00000;
22177 : 00000;
22200 : 00000;
22201 : 00000;
22202 : 00000;
22203 : 00000;
22204 : 00000;
22205 : 00000;
22206 : 00000;
22207 : 00000;
22210 : 00000;
22211 : 00000;
22212 : 00000;
22213 : 00000;
22214 : 00000;
22215 : 00000;
22216 : 00000;
22217 : 00000;
22220 : 00000;
22221 : 00000;
22222 : 00000;
22223 : 00000;
22224 : 00000;
22225 : 00000;
22226 : 00000;
22227 : 00000;
22230 : 00000;
22231 : 00000;
22232 : 00000;
22233 : 00000;
22234 : 00000;
22235 : 00000;
22236 : 00000;
22237 : 00000;
22240 : 00000;
22241 : 00000;
22242 : 00000;
22243 : 00000;
22244 : 00000;
22245 : 00000;
22246 : 00000;
22247 : 00000;
22250 : 00000;
22251 : 00000;
22252 : 00000;
22253 : 00000;
22254 : 00000;
22255 : 00000;
22256 : 00000;
22257 : 00000;
22260 : 00000;
22261 : 00000;
22262 : 00000;
22263 : 00000;
22264 : 00000;
22265 : 00000;
22266 : 00000;
22267 : 00000;
22270 : 00000;
22271 : 00000;
22272 : 00000;
22273 : 00000;
22274 : 00000;
22275 : 00000;
22276 : 00000;
22277 : 00000;
22300 : 00000;
22301 : 00000;
22302 : 00000;
22303 : 00000;
22304 : 00000;
22305 : 00000;
22306 : 00000;
22307 : 00000;
22310 : 00000;
22311 : 00000;
22312 : 00000;
22313 : 00000;
22314 : 00000;
22315 : 00000;
22316 : 00000;
22317 : 00000;
22320 : 00000;
22321 : 00000;
22322 : 00000;
22323 : 00000;
22324 : 00000;
22325 : 00000;
22326 : 00000;
22327 : 00000;
22330 : 00000;
22331 : 00000;
22332 : 00000;
22333 : 00000;
22334 : 00000;
22335 : 00000;
22336 : 00000;
22337 : 00000;
22340 : 00000;
22341 : 00000;
22342 : 00000;
22343 : 00000;
22344 : 00000;
22345 : 00000;
22346 : 00000;
22347 : 00000;
22350 : 00000;
22351 : 00000;
22352 : 00000;
22353 : 00000;
22354 : 00000;
22355 : 00000;
22356 : 00000;
22357 : 00000;
22360 : 00000;
22361 : 00000;
22362 : 00000;
22363 : 00000;
22364 : 00000;
22365 : 00000;
22366 : 00000;
22367 : 00000;
22370 : 00000;
22371 : 00000;
22372 : 00000;
22373 : 00000;
22374 : 00000;
22375 : 00000;
22376 : 00000;
22377 : 00000;
22400 : 00000;
22401 : 00000;
22402 : 00000;
22403 : 00000;
22404 : 00000;
22405 : 00000;
22406 : 00000;
22407 : 00000;
22410 : 00000;
22411 : 00000;
22412 : 00000;
22413 : 00000;
22414 : 00000;
22415 : 00000;
22416 : 00000;
22417 : 00000;
22420 : 00000;
22421 : 00000;
22422 : 00000;
22423 : 00000;
22424 : 00000;
22425 : 00000;
22426 : 00000;
22427 : 00000;
22430 : 00000;
22431 : 00000;
22432 : 00000;
22433 : 00000;
22434 : 00000;
22435 : 00000;
22436 : 00000;
22437 : 00000;
22440 : 00000;
22441 : 00000;
22442 : 00000;
22443 : 00000;
22444 : 00000;
22445 : 00000;
22446 : 00000;
22447 : 00000;
22450 : 00000;
22451 : 00000;
22452 : 00000;
22453 : 00000;
22454 : 00000;
22455 : 00000;
22456 : 00000;
22457 : 00000;
22460 : 00000;
22461 : 00000;
22462 : 00000;
22463 : 00000;
22464 : 00000;
22465 : 00000;
22466 : 00000;
22467 : 00000;
22470 : 00000;
22471 : 00000;
22472 : 00000;
22473 : 00000;
22474 : 00000;
22475 : 00000;
22476 : 00000;
22477 : 00000;
22500 : 00000;
22501 : 00000;
22502 : 00000;
22503 : 00000;
22504 : 00000;
22505 : 00000;
22506 : 00000;
22507 : 00000;
22510 : 00000;
22511 : 00000;
22512 : 00000;
22513 : 00000;
22514 : 00000;
22515 : 00000;
22516 : 00000;
22517 : 00000;
22520 : 00000;
22521 : 00000;
22522 : 00000;
22523 : 00000;
22524 : 00000;
22525 : 00000;
22526 : 00000;
22527 : 00000;
22530 : 00000;
22531 : 00000;
22532 : 00000;
22533 : 00000;
22534 : 00000;
22535 : 00000;
22536 : 00000;
22537 : 00000;
22540 : 00000;
22541 : 00000;
22542 : 00000;
22543 : 00000;
22544 : 00000;
22545 : 00000;
22546 : 00000;
22547 : 00000;
22550 : 00000;
22551 : 00000;
22552 : 00000;
22553 : 00000;
22554 : 00000;
22555 : 00000;
22556 : 00000;
22557 : 00000;
22560 : 00000;
22561 : 00000;
22562 : 00000;
22563 : 00000;
22564 : 00000;
22565 : 00000;
22566 : 00000;
22567 : 00000;
22570 : 00000;
22571 : 00000;
22572 : 00000;
22573 : 00000;
22574 : 00000;
22575 : 00000;
22576 : 00000;
22577 : 00000;
22600 : 00000;
22601 : 00000;
22602 : 00000;
22603 : 00000;
22604 : 00000;
22605 : 00000;
22606 : 00000;
22607 : 00000;
22610 : 00000;
22611 : 00000;
22612 : 00000;
22613 : 00000;
22614 : 00000;
22615 : 00000;
22616 : 00000;
22617 : 00000;
22620 : 00000;
22621 : 00000;
22622 : 00000;
22623 : 00000;
22624 : 00000;
22625 : 00000;
22626 : 00000;
22627 : 00000;
22630 : 00000;
22631 : 00000;
22632 : 00000;
22633 : 00000;
22634 : 00000;
22635 : 00000;
22636 : 00000;
22637 : 00000;
22640 : 00000;
22641 : 00000;
22642 : 00000;
22643 : 00000;
22644 : 00000;
22645 : 00000;
22646 : 00000;
22647 : 00000;
22650 : 00000;
22651 : 00000;
22652 : 00000;
22653 : 00000;
22654 : 00000;
22655 : 00000;
22656 : 00000;
22657 : 00000;
22660 : 00000;
22661 : 00000;
22662 : 00000;
22663 : 00000;
22664 : 00000;
22665 : 00000;
22666 : 00000;
22667 : 00000;
22670 : 00000;
22671 : 00000;
22672 : 00000;
22673 : 00000;
22674 : 00000;
22675 : 00000;
22676 : 00000;
22677 : 00000;
22700 : 00000;
22701 : 00000;
22702 : 00000;
22703 : 00000;
22704 : 00000;
22705 : 00000;
22706 : 00000;
22707 : 00000;
22710 : 00000;
22711 : 00000;
22712 : 00000;
22713 : 00000;
22714 : 00000;
22715 : 00000;
22716 : 00000;
22717 : 00000;
22720 : 00000;
22721 : 00000;
22722 : 00000;
22723 : 00000;
22724 : 00000;
22725 : 00000;
22726 : 00000;
22727 : 00000;
22730 : 00000;
22731 : 00000;
22732 : 00000;
22733 : 00000;
22734 : 00000;
22735 : 00000;
22736 : 00000;
22737 : 00000;
22740 : 00000;
22741 : 00000;
22742 : 00000;
22743 : 00000;
22744 : 00000;
22745 : 00000;
22746 : 00000;
22747 : 00000;
22750 : 00000;
22751 : 00000;
22752 : 00000;
22753 : 00000;
22754 : 00000;
22755 : 00000;
22756 : 00000;
22757 : 00000;
22760 : 00000;
22761 : 00000;
22762 : 00000;
22763 : 00000;
22764 : 00000;
22765 : 00000;
22766 : 00000;
22767 : 00000;
22770 : 00000;
22771 : 00000;
22772 : 00000;
22773 : 00000;
22774 : 00000;
22775 : 00000;
22776 : 00000;
22777 : 00000;
23000 : 00000;
23001 : 00000;
23002 : 00000;
23003 : 00000;
23004 : 00000;
23005 : 00000;
23006 : 00000;
23007 : 00000;
23010 : 00000;
23011 : 00000;
23012 : 00000;
23013 : 00000;
23014 : 00000;
23015 : 00000;
23016 : 00000;
23017 : 00000;
23020 : 00000;
23021 : 00000;
23022 : 00000;
23023 : 00000;
23024 : 00000;
23025 : 00000;
23026 : 00000;
23027 : 00000;
23030 : 00000;
23031 : 00000;
23032 : 00000;
23033 : 00000;
23034 : 00000;
23035 : 00000;
23036 : 00000;
23037 : 00000;
23040 : 00000;
23041 : 00000;
23042 : 00000;
23043 : 00000;
23044 : 00000;
23045 : 00000;
23046 : 00000;
23047 : 00000;
23050 : 00000;
23051 : 00000;
23052 : 00000;
23053 : 00000;
23054 : 00000;
23055 : 00000;
23056 : 00000;
23057 : 00000;
23060 : 00000;
23061 : 00000;
23062 : 00000;
23063 : 00000;
23064 : 00000;
23065 : 00000;
23066 : 00000;
23067 : 00000;
23070 : 00000;
23071 : 00000;
23072 : 00000;
23073 : 00000;
23074 : 00000;
23075 : 00000;
23076 : 00000;
23077 : 00000;
23100 : 00000;
23101 : 00000;
23102 : 00000;
23103 : 00000;
23104 : 00000;
23105 : 00000;
23106 : 00000;
23107 : 00000;
23110 : 00000;
23111 : 00000;
23112 : 00000;
23113 : 00000;
23114 : 00000;
23115 : 00000;
23116 : 00000;
23117 : 00000;
23120 : 00000;
23121 : 00000;
23122 : 00000;
23123 : 00000;
23124 : 00000;
23125 : 00000;
23126 : 00000;
23127 : 00000;
23130 : 00000;
23131 : 00000;
23132 : 00000;
23133 : 00000;
23134 : 00000;
23135 : 00000;
23136 : 00000;
23137 : 00000;
23140 : 00000;
23141 : 00000;
23142 : 00000;
23143 : 00000;
23144 : 00000;
23145 : 00000;
23146 : 00000;
23147 : 00000;
23150 : 00000;
23151 : 00000;
23152 : 00000;
23153 : 00000;
23154 : 00000;
23155 : 00000;
23156 : 00000;
23157 : 00000;
23160 : 00000;
23161 : 00000;
23162 : 00000;
23163 : 00000;
23164 : 00000;
23165 : 00000;
23166 : 00000;
23167 : 00000;
23170 : 00000;
23171 : 00000;
23172 : 00000;
23173 : 00000;
23174 : 00000;
23175 : 00000;
23176 : 00000;
23177 : 00000;
23200 : 00000;
23201 : 00000;
23202 : 00000;
23203 : 00000;
23204 : 00000;
23205 : 00000;
23206 : 00000;
23207 : 00000;
23210 : 00000;
23211 : 00000;
23212 : 00000;
23213 : 00000;
23214 : 00000;
23215 : 00000;
23216 : 00000;
23217 : 00000;
23220 : 00000;
23221 : 00000;
23222 : 00000;
23223 : 00000;
23224 : 00000;
23225 : 00000;
23226 : 00000;
23227 : 00000;
23230 : 00000;
23231 : 00000;
23232 : 00000;
23233 : 00000;
23234 : 00000;
23235 : 00000;
23236 : 00000;
23237 : 00000;
23240 : 00000;
23241 : 00000;
23242 : 00000;
23243 : 00000;
23244 : 00000;
23245 : 00000;
23246 : 00000;
23247 : 00000;
23250 : 00000;
23251 : 00000;
23252 : 00000;
23253 : 00000;
23254 : 00000;
23255 : 00000;
23256 : 00000;
23257 : 00000;
23260 : 00000;
23261 : 00000;
23262 : 00000;
23263 : 00000;
23264 : 00000;
23265 : 00000;
23266 : 00000;
23267 : 00000;
23270 : 00000;
23271 : 00000;
23272 : 00000;
23273 : 00000;
23274 : 00000;
23275 : 00000;
23276 : 00000;
23277 : 00000;
23300 : 00000;
23301 : 00000;
23302 : 00000;
23303 : 00000;
23304 : 00000;
23305 : 00000;
23306 : 00000;
23307 : 00000;
23310 : 00000;
23311 : 00000;
23312 : 00000;
23313 : 00000;
23314 : 00000;
23315 : 00000;
23316 : 00000;
23317 : 00000;
23320 : 00000;
23321 : 00000;
23322 : 00000;
23323 : 00000;
23324 : 00000;
23325 : 00000;
23326 : 00000;
23327 : 00000;
23330 : 00000;
23331 : 00000;
23332 : 00000;
23333 : 00000;
23334 : 00000;
23335 : 00000;
23336 : 00000;
23337 : 00000;
23340 : 00000;
23341 : 00000;
23342 : 00000;
23343 : 00000;
23344 : 00000;
23345 : 00000;
23346 : 00000;
23347 : 00000;
23350 : 00000;
23351 : 00000;
23352 : 00000;
23353 : 00000;
23354 : 00000;
23355 : 00000;
23356 : 00000;
23357 : 00000;
23360 : 00000;
23361 : 00000;
23362 : 00000;
23363 : 00000;
23364 : 00000;
23365 : 00000;
23366 : 00000;
23367 : 00000;
23370 : 00000;
23371 : 00000;
23372 : 00000;
23373 : 00000;
23374 : 00000;
23375 : 00000;
23376 : 00000;
23377 : 00000;
23400 : 00000;
23401 : 00000;
23402 : 00000;
23403 : 00000;
23404 : 00000;
23405 : 00000;
23406 : 00000;
23407 : 00000;
23410 : 00000;
23411 : 00000;
23412 : 00000;
23413 : 00000;
23414 : 00000;
23415 : 00000;
23416 : 00000;
23417 : 00000;
23420 : 00000;
23421 : 00000;
23422 : 00000;
23423 : 00000;
23424 : 00000;
23425 : 00000;
23426 : 00000;
23427 : 00000;
23430 : 00000;
23431 : 00000;
23432 : 00000;
23433 : 00000;
23434 : 00000;
23435 : 00000;
23436 : 00000;
23437 : 00000;
23440 : 00000;
23441 : 00000;
23442 : 00000;
23443 : 00000;
23444 : 00000;
23445 : 00000;
23446 : 00000;
23447 : 00000;
23450 : 00000;
23451 : 00000;
23452 : 00000;
23453 : 00000;
23454 : 00000;
23455 : 00000;
23456 : 00000;
23457 : 00000;
23460 : 00000;
23461 : 00000;
23462 : 00000;
23463 : 00000;
23464 : 00000;
23465 : 00000;
23466 : 00000;
23467 : 00000;
23470 : 00000;
23471 : 00000;
23472 : 00000;
23473 : 00000;
23474 : 00000;
23475 : 00000;
23476 : 00000;
23477 : 00000;
23500 : 00000;
23501 : 00000;
23502 : 00000;
23503 : 00000;
23504 : 00000;
23505 : 00000;
23506 : 00000;
23507 : 00000;
23510 : 00000;
23511 : 00000;
23512 : 00000;
23513 : 00000;
23514 : 00000;
23515 : 00000;
23516 : 00000;
23517 : 00000;
23520 : 00000;
23521 : 00000;
23522 : 00000;
23523 : 00000;
23524 : 00000;
23525 : 00000;
23526 : 00000;
23527 : 00000;
23530 : 00000;
23531 : 00000;
23532 : 00000;
23533 : 00000;
23534 : 00000;
23535 : 00000;
23536 : 00000;
23537 : 00000;
23540 : 00000;
23541 : 00000;
23542 : 00000;
23543 : 00000;
23544 : 00000;
23545 : 00000;
23546 : 00000;
23547 : 00000;
23550 : 00000;
23551 : 00000;
23552 : 00000;
23553 : 00000;
23554 : 00000;
23555 : 00000;
23556 : 00000;
23557 : 00000;
23560 : 00000;
23561 : 00000;
23562 : 00000;
23563 : 00000;
23564 : 00000;
23565 : 00000;
23566 : 00000;
23567 : 00000;
23570 : 00000;
23571 : 00000;
23572 : 00000;
23573 : 00000;
23574 : 00000;
23575 : 00000;
23576 : 00000;
23577 : 00000;
23600 : 00000;
23601 : 00000;
23602 : 00000;
23603 : 00000;
23604 : 00000;
23605 : 00000;
23606 : 00000;
23607 : 00000;
23610 : 00000;
23611 : 00000;
23612 : 00000;
23613 : 00000;
23614 : 00000;
23615 : 00000;
23616 : 00000;
23617 : 00000;
23620 : 00000;
23621 : 00000;
23622 : 00000;
23623 : 00000;
23624 : 00000;
23625 : 00000;
23626 : 00000;
23627 : 00000;
23630 : 00000;
23631 : 00000;
23632 : 00000;
23633 : 00000;
23634 : 00000;
23635 : 00000;
23636 : 00000;
23637 : 00000;
23640 : 00000;
23641 : 00000;
23642 : 00000;
23643 : 00000;
23644 : 00000;
23645 : 00000;
23646 : 00000;
23647 : 00000;
23650 : 00000;
23651 : 00000;
23652 : 00000;
23653 : 00000;
23654 : 00000;
23655 : 00000;
23656 : 00000;
23657 : 00000;
23660 : 00000;
23661 : 00000;
23662 : 00000;
23663 : 00000;
23664 : 00000;
23665 : 00000;
23666 : 00000;
23667 : 00000;
23670 : 00000;
23671 : 00000;
23672 : 00000;
23673 : 00000;
23674 : 00000;
23675 : 00000;
23676 : 00000;
23677 : 00000;
23700 : 00000;
23701 : 00000;
23702 : 00000;
23703 : 00000;
23704 : 00000;
23705 : 00000;
23706 : 00000;
23707 : 00000;
23710 : 00000;
23711 : 00000;
23712 : 00000;
23713 : 00000;
23714 : 00000;
23715 : 00000;
23716 : 00000;
23717 : 00000;
23720 : 00000;
23721 : 00000;
23722 : 00000;
23723 : 00000;
23724 : 00000;
23725 : 00000;
23726 : 00000;
23727 : 00000;
23730 : 00000;
23731 : 00000;
23732 : 00000;
23733 : 00000;
23734 : 00000;
23735 : 00000;
23736 : 00000;
23737 : 00000;
23740 : 00000;
23741 : 00000;
23742 : 00000;
23743 : 00000;
23744 : 00000;
23745 : 00000;
23746 : 00000;
23747 : 00000;
23750 : 00000;
23751 : 00000;
23752 : 00000;
23753 : 00000;
23754 : 00000;
23755 : 00000;
23756 : 00000;
23757 : 00000;
23760 : 00000;
23761 : 00000;
23762 : 00000;
23763 : 00000;
23764 : 00000;
23765 : 00000;
23766 : 00000;
23767 : 00000;
23770 : 00000;
23771 : 00000;
23772 : 00000;
23773 : 00000;
23774 : 00000;
23775 : 00000;
23776 : 00000;
23777 : 00000;
24000 : 00000;
24001 : 00000;
24002 : 00000;
24003 : 00000;
24004 : 00000;
24005 : 00000;
24006 : 00000;
24007 : 00000;
24010 : 00000;
24011 : 00000;
24012 : 00000;
24013 : 00000;
24014 : 00000;
24015 : 00000;
24016 : 00000;
24017 : 00000;
24020 : 00000;
24021 : 00000;
24022 : 00000;
24023 : 00000;
24024 : 00000;
24025 : 00000;
24026 : 00000;
24027 : 00000;
24030 : 00000;
24031 : 00000;
24032 : 00000;
24033 : 00000;
24034 : 00000;
24035 : 00000;
24036 : 00000;
24037 : 00000;
24040 : 00000;
24041 : 00000;
24042 : 00000;
24043 : 00000;
24044 : 00000;
24045 : 00000;
24046 : 00000;
24047 : 00000;
24050 : 00000;
24051 : 00000;
24052 : 00000;
24053 : 00000;
24054 : 00000;
24055 : 00000;
24056 : 00000;
24057 : 00000;
24060 : 00000;
24061 : 00000;
24062 : 00000;
24063 : 00000;
24064 : 00000;
24065 : 00000;
24066 : 00000;
24067 : 00000;
24070 : 00000;
24071 : 00000;
24072 : 00000;
24073 : 00000;
24074 : 00000;
24075 : 00000;
24076 : 00000;
24077 : 00000;
24100 : 00000;
24101 : 00000;
24102 : 00000;
24103 : 00000;
24104 : 00000;
24105 : 00000;
24106 : 00000;
24107 : 00000;
24110 : 00000;
24111 : 00000;
24112 : 00000;
24113 : 00000;
24114 : 00000;
24115 : 00000;
24116 : 00000;
24117 : 00000;
24120 : 00000;
24121 : 00000;
24122 : 00000;
24123 : 00000;
24124 : 00000;
24125 : 00000;
24126 : 00000;
24127 : 00000;
24130 : 00000;
24131 : 00000;
24132 : 00000;
24133 : 00000;
24134 : 00000;
24135 : 00000;
24136 : 00000;
24137 : 00000;
24140 : 00000;
24141 : 00000;
24142 : 00000;
24143 : 00000;
24144 : 00000;
24145 : 00000;
24146 : 00000;
24147 : 00000;
24150 : 00000;
24151 : 00000;
24152 : 00000;
24153 : 00000;
24154 : 00000;
24155 : 00000;
24156 : 00000;
24157 : 00000;
24160 : 00000;
24161 : 00000;
24162 : 00000;
24163 : 00000;
24164 : 00000;
24165 : 00000;
24166 : 00000;
24167 : 00000;
24170 : 00000;
24171 : 00000;
24172 : 00000;
24173 : 00000;
24174 : 00000;
24175 : 00000;
24176 : 00000;
24177 : 00000;
24200 : 00000;
24201 : 00000;
24202 : 00000;
24203 : 00000;
24204 : 00000;
24205 : 00000;
24206 : 00000;
24207 : 00000;
24210 : 00000;
24211 : 00000;
24212 : 00000;
24213 : 00000;
24214 : 00000;
24215 : 00000;
24216 : 00000;
24217 : 00000;
24220 : 00000;
24221 : 00000;
24222 : 00000;
24223 : 00000;
24224 : 00000;
24225 : 00000;
24226 : 00000;
24227 : 00000;
24230 : 00000;
24231 : 00000;
24232 : 00000;
24233 : 00000;
24234 : 00000;
24235 : 00000;
24236 : 00000;
24237 : 00000;
24240 : 00000;
24241 : 00000;
24242 : 00000;
24243 : 00000;
24244 : 00000;
24245 : 00000;
24246 : 00000;
24247 : 00000;
24250 : 00000;
24251 : 00000;
24252 : 00000;
24253 : 00000;
24254 : 00000;
24255 : 00000;
24256 : 00000;
24257 : 00000;
24260 : 00000;
24261 : 00000;
24262 : 00000;
24263 : 00000;
24264 : 00000;
24265 : 00000;
24266 : 00000;
24267 : 00000;
24270 : 00000;
24271 : 00000;
24272 : 00000;
24273 : 00000;
24274 : 00000;
24275 : 00000;
24276 : 00000;
24277 : 00000;
24300 : 00000;
24301 : 00000;
24302 : 00000;
24303 : 00000;
24304 : 00000;
24305 : 00000;
24306 : 00000;
24307 : 00000;
24310 : 00000;
24311 : 00000;
24312 : 00000;
24313 : 00000;
24314 : 00000;
24315 : 00000;
24316 : 00000;
24317 : 00000;
24320 : 00000;
24321 : 00000;
24322 : 00000;
24323 : 00000;
24324 : 00000;
24325 : 00000;
24326 : 00000;
24327 : 00000;
24330 : 00000;
24331 : 00000;
24332 : 00000;
24333 : 00000;
24334 : 00000;
24335 : 00000;
24336 : 00000;
24337 : 00000;
24340 : 00000;
24341 : 00000;
24342 : 00000;
24343 : 00000;
24344 : 00000;
24345 : 00000;
24346 : 00000;
24347 : 00000;
24350 : 00000;
24351 : 00000;
24352 : 00000;
24353 : 00000;
24354 : 00000;
24355 : 00000;
24356 : 00000;
24357 : 00000;
24360 : 00000;
24361 : 00000;
24362 : 00000;
24363 : 00000;
24364 : 00000;
24365 : 00000;
24366 : 00000;
24367 : 00000;
24370 : 00000;
24371 : 00000;
24372 : 00000;
24373 : 00000;
24374 : 00000;
24375 : 00000;
24376 : 00000;
24377 : 00000;
24400 : 00000;
24401 : 00000;
24402 : 00000;
24403 : 00000;
24404 : 00000;
24405 : 00000;
24406 : 00000;
24407 : 00000;
24410 : 00000;
24411 : 00000;
24412 : 00000;
24413 : 00000;
24414 : 00000;
24415 : 00000;
24416 : 00000;
24417 : 00000;
24420 : 00000;
24421 : 00000;
24422 : 00000;
24423 : 00000;
24424 : 00000;
24425 : 00000;
24426 : 00000;
24427 : 00000;
24430 : 00000;
24431 : 00000;
24432 : 00000;
24433 : 00000;
24434 : 00000;
24435 : 00000;
24436 : 00000;
24437 : 00000;
24440 : 00000;
24441 : 00000;
24442 : 00000;
24443 : 00000;
24444 : 00000;
24445 : 00000;
24446 : 00000;
24447 : 00000;
24450 : 00000;
24451 : 00000;
24452 : 00000;
24453 : 00000;
24454 : 00000;
24455 : 00000;
24456 : 00000;
24457 : 00000;
24460 : 00000;
24461 : 00000;
24462 : 00000;
24463 : 00000;
24464 : 00000;
24465 : 00000;
24466 : 00000;
24467 : 00000;
24470 : 00000;
24471 : 00000;
24472 : 00000;
24473 : 00000;
24474 : 00000;
24475 : 00000;
24476 : 00000;
24477 : 00000;
24500 : 00000;
24501 : 00000;
24502 : 00000;
24503 : 00000;
24504 : 00000;
24505 : 00000;
24506 : 00000;
24507 : 00000;
24510 : 00000;
24511 : 00000;
24512 : 00000;
24513 : 00000;
24514 : 00000;
24515 : 00000;
24516 : 00000;
24517 : 00000;
24520 : 00000;
24521 : 00000;
24522 : 00000;
24523 : 00000;
24524 : 00000;
24525 : 00000;
24526 : 00000;
24527 : 00000;
24530 : 00000;
24531 : 00000;
24532 : 00000;
24533 : 00000;
24534 : 00000;
24535 : 00000;
24536 : 00000;
24537 : 00000;
24540 : 00000;
24541 : 00000;
24542 : 00000;
24543 : 00000;
24544 : 00000;
24545 : 00000;
24546 : 00000;
24547 : 00000;
24550 : 00000;
24551 : 00000;
24552 : 00000;
24553 : 00000;
24554 : 00000;
24555 : 00000;
24556 : 00000;
24557 : 00000;
24560 : 00000;
24561 : 00000;
24562 : 00000;
24563 : 00000;
24564 : 00000;
24565 : 00000;
24566 : 00000;
24567 : 00000;
24570 : 00000;
24571 : 00000;
24572 : 00000;
24573 : 00000;
24574 : 00000;
24575 : 00000;
24576 : 00000;
24577 : 00000;
24600 : 00000;
24601 : 00000;
24602 : 00000;
24603 : 00000;
24604 : 00000;
24605 : 00000;
24606 : 00000;
24607 : 00000;
24610 : 00000;
24611 : 00000;
24612 : 00000;
24613 : 00000;
24614 : 00000;
24615 : 00000;
24616 : 00000;
24617 : 00000;
24620 : 00000;
24621 : 00000;
24622 : 00000;
24623 : 00000;
24624 : 00000;
24625 : 00000;
24626 : 00000;
24627 : 00000;
24630 : 00000;
24631 : 00000;
24632 : 00000;
24633 : 00000;
24634 : 00000;
24635 : 00000;
24636 : 00000;
24637 : 00000;
24640 : 00000;
24641 : 00000;
24642 : 00000;
24643 : 00000;
24644 : 00000;
24645 : 00000;
24646 : 00000;
24647 : 00000;
24650 : 00000;
24651 : 00000;
24652 : 00000;
24653 : 00000;
24654 : 00000;
24655 : 00000;
24656 : 00000;
24657 : 00000;
24660 : 00000;
24661 : 00000;
24662 : 00000;
24663 : 00000;
24664 : 00000;
24665 : 00000;
24666 : 00000;
24667 : 00000;
24670 : 00000;
24671 : 00000;
24672 : 00000;
24673 : 00000;
24674 : 00000;
24675 : 00000;
24676 : 00000;
24677 : 00000;
24700 : 00000;
24701 : 00000;
24702 : 00000;
24703 : 00000;
24704 : 00000;
24705 : 00000;
24706 : 00000;
24707 : 00000;
24710 : 00000;
24711 : 00000;
24712 : 00000;
24713 : 00000;
24714 : 00000;
24715 : 00000;
24716 : 00000;
24717 : 00000;
24720 : 00000;
24721 : 00000;
24722 : 00000;
24723 : 00000;
24724 : 00000;
24725 : 00000;
24726 : 00000;
24727 : 00000;
24730 : 00000;
24731 : 00000;
24732 : 00000;
24733 : 00000;
24734 : 00000;
24735 : 00000;
24736 : 00000;
24737 : 00000;
24740 : 00000;
24741 : 00000;
24742 : 00000;
24743 : 00000;
24744 : 00000;
24745 : 00000;
24746 : 00000;
24747 : 00000;
24750 : 00000;
24751 : 00000;
24752 : 00000;
24753 : 00000;
24754 : 00000;
24755 : 00000;
24756 : 00000;
24757 : 00000;
24760 : 00000;
24761 : 00000;
24762 : 00000;
24763 : 00000;
24764 : 00000;
24765 : 00000;
24766 : 00000;
24767 : 00000;
24770 : 00000;
24771 : 00000;
24772 : 00000;
24773 : 00000;
24774 : 00000;
24775 : 00000;
24776 : 00000;
24777 : 00000;
25000 : 00000;
25001 : 00000;
25002 : 00000;
25003 : 00000;
25004 : 00000;
25005 : 00000;
25006 : 00000;
25007 : 00000;
25010 : 00000;
25011 : 00000;
25012 : 00000;
25013 : 00000;
25014 : 00000;
25015 : 00000;
25016 : 00000;
25017 : 00000;
25020 : 00000;
25021 : 00000;
25022 : 00000;
25023 : 00000;
25024 : 00000;
25025 : 00000;
25026 : 00000;
25027 : 00000;
25030 : 00000;
25031 : 00000;
25032 : 00000;
25033 : 00000;
25034 : 00000;
25035 : 00000;
25036 : 00000;
25037 : 00000;
25040 : 00000;
25041 : 00000;
25042 : 00000;
25043 : 00000;
25044 : 00000;
25045 : 00000;
25046 : 00000;
25047 : 00000;
25050 : 00000;
25051 : 00000;
25052 : 00000;
25053 : 00000;
25054 : 00000;
25055 : 00000;
25056 : 00000;
25057 : 00000;
25060 : 00000;
25061 : 00000;
25062 : 00000;
25063 : 00000;
25064 : 00000;
25065 : 00000;
25066 : 00000;
25067 : 00000;
25070 : 00000;
25071 : 00000;
25072 : 00000;
25073 : 00000;
25074 : 00000;
25075 : 00000;
25076 : 00000;
25077 : 00000;
25100 : 00000;
25101 : 00000;
25102 : 00000;
25103 : 00000;
25104 : 00000;
25105 : 00000;
25106 : 00000;
25107 : 00000;
25110 : 00000;
25111 : 00000;
25112 : 00000;
25113 : 00000;
25114 : 00000;
25115 : 00000;
25116 : 00000;
25117 : 00000;
25120 : 00000;
25121 : 00000;
25122 : 00000;
25123 : 00000;
25124 : 00000;
25125 : 00000;
25126 : 00000;
25127 : 00000;
25130 : 00000;
25131 : 00000;
25132 : 00000;
25133 : 00000;
25134 : 00000;
25135 : 00000;
25136 : 00000;
25137 : 00000;
25140 : 00000;
25141 : 00000;
25142 : 00000;
25143 : 00000;
25144 : 00000;
25145 : 00000;
25146 : 00000;
25147 : 00000;
25150 : 00000;
25151 : 00000;
25152 : 00000;
25153 : 00000;
25154 : 00000;
25155 : 00000;
25156 : 00000;
25157 : 00000;
25160 : 00000;
25161 : 00000;
25162 : 00000;
25163 : 00000;
25164 : 00000;
25165 : 00000;
25166 : 00000;
25167 : 00000;
25170 : 00000;
25171 : 00000;
25172 : 00000;
25173 : 00000;
25174 : 00000;
25175 : 00000;
25176 : 00000;
25177 : 00000;
25200 : 00000;
25201 : 00000;
25202 : 00000;
25203 : 00000;
25204 : 00000;
25205 : 00000;
25206 : 00000;
25207 : 00000;
25210 : 00000;
25211 : 00000;
25212 : 00000;
25213 : 00000;
25214 : 00000;
25215 : 00000;
25216 : 00000;
25217 : 00000;
25220 : 00000;
25221 : 00000;
25222 : 00000;
25223 : 00000;
25224 : 00000;
25225 : 00000;
25226 : 00000;
25227 : 00000;
25230 : 00000;
25231 : 00000;
25232 : 00000;
25233 : 00000;
25234 : 00000;
25235 : 00000;
25236 : 00000;
25237 : 00000;
25240 : 00000;
25241 : 00000;
25242 : 00000;
25243 : 00000;
25244 : 00000;
25245 : 00000;
25246 : 00000;
25247 : 00000;
25250 : 00000;
25251 : 00000;
25252 : 00000;
25253 : 00000;
25254 : 00000;
25255 : 00000;
25256 : 00000;
25257 : 00000;
25260 : 00000;
25261 : 00000;
25262 : 00000;
25263 : 00000;
25264 : 00000;
25265 : 00000;
25266 : 00000;
25267 : 00000;
25270 : 00000;
25271 : 00000;
25272 : 00000;
25273 : 00000;
25274 : 00000;
25275 : 00000;
25276 : 00000;
25277 : 00000;
25300 : 00000;
25301 : 00000;
25302 : 00000;
25303 : 00000;
25304 : 00000;
25305 : 00000;
25306 : 00000;
25307 : 00000;
25310 : 00000;
25311 : 00000;
25312 : 00000;
25313 : 00000;
25314 : 00000;
25315 : 00000;
25316 : 00000;
25317 : 00000;
25320 : 00000;
25321 : 00000;
25322 : 00000;
25323 : 00000;
25324 : 00000;
25325 : 00000;
25326 : 00000;
25327 : 00000;
25330 : 00000;
25331 : 00000;
25332 : 00000;
25333 : 00000;
25334 : 00000;
25335 : 00000;
25336 : 00000;
25337 : 00000;
25340 : 00000;
25341 : 00000;
25342 : 00000;
25343 : 00000;
25344 : 00000;
25345 : 00000;
25346 : 00000;
25347 : 00000;
25350 : 00000;
25351 : 00000;
25352 : 00000;
25353 : 00000;
25354 : 00000;
25355 : 00000;
25356 : 00000;
25357 : 00000;
25360 : 00000;
25361 : 00000;
25362 : 00000;
25363 : 00000;
25364 : 00000;
25365 : 00000;
25366 : 00000;
25367 : 00000;
25370 : 00000;
25371 : 00000;
25372 : 00000;
25373 : 00000;
25374 : 00000;
25375 : 00000;
25376 : 00000;
25377 : 00000;
25400 : 00000;
25401 : 00000;
25402 : 00000;
25403 : 00000;
25404 : 00000;
25405 : 00000;
25406 : 00000;
25407 : 00000;
25410 : 00000;
25411 : 00000;
25412 : 00000;
25413 : 00000;
25414 : 00000;
25415 : 00000;
25416 : 00000;
25417 : 00000;
25420 : 00000;
25421 : 00000;
25422 : 00000;
25423 : 00000;
25424 : 00000;
25425 : 00000;
25426 : 00000;
25427 : 00000;
25430 : 00000;
25431 : 00000;
25432 : 00000;
25433 : 00000;
25434 : 00000;
25435 : 00000;
25436 : 00000;
25437 : 00000;
25440 : 00000;
25441 : 00000;
25442 : 00000;
25443 : 00000;
25444 : 00000;
25445 : 00000;
25446 : 00000;
25447 : 00000;
25450 : 00000;
25451 : 00000;
25452 : 00000;
25453 : 00000;
25454 : 00000;
25455 : 00000;
25456 : 00000;
25457 : 00000;
25460 : 00000;
25461 : 00000;
25462 : 00000;
25463 : 00000;
25464 : 00000;
25465 : 00000;
25466 : 00000;
25467 : 00000;
25470 : 00000;
25471 : 00000;
25472 : 00000;
25473 : 00000;
25474 : 00000;
25475 : 00000;
25476 : 00000;
25477 : 00000;
25500 : 00000;
25501 : 00000;
25502 : 00000;
25503 : 00000;
25504 : 00000;
25505 : 00000;
25506 : 00000;
25507 : 00000;
25510 : 00000;
25511 : 00000;
25512 : 00000;
25513 : 00000;
25514 : 00000;
25515 : 00000;
25516 : 00000;
25517 : 00000;
25520 : 00000;
25521 : 00000;
25522 : 00000;
25523 : 00000;
25524 : 00000;
25525 : 00000;
25526 : 00000;
25527 : 00000;
25530 : 00000;
25531 : 00000;
25532 : 00000;
25533 : 00000;
25534 : 00000;
25535 : 00000;
25536 : 00000;
25537 : 00000;
25540 : 00000;
25541 : 00000;
25542 : 00000;
25543 : 00000;
25544 : 00000;
25545 : 00000;
25546 : 00000;
25547 : 00000;
25550 : 00000;
25551 : 00000;
25552 : 00000;
25553 : 00000;
25554 : 00000;
25555 : 00000;
25556 : 00000;
25557 : 00000;
25560 : 00000;
25561 : 00000;
25562 : 00000;
25563 : 00000;
25564 : 00000;
25565 : 00000;
25566 : 00000;
25567 : 00000;
25570 : 00000;
25571 : 00000;
25572 : 00000;
25573 : 00000;
25574 : 00000;
25575 : 00000;
25576 : 00000;
25577 : 00000;
25600 : 00000;
25601 : 00000;
25602 : 00000;
25603 : 00000;
25604 : 00000;
25605 : 00000;
25606 : 00000;
25607 : 00000;
25610 : 00000;
25611 : 00000;
25612 : 00000;
25613 : 00000;
25614 : 00000;
25615 : 00000;
25616 : 00000;
25617 : 00000;
25620 : 00000;
25621 : 00000;
25622 : 00000;
25623 : 00000;
25624 : 00000;
25625 : 00000;
25626 : 00000;
25627 : 00000;
25630 : 00000;
25631 : 00000;
25632 : 00000;
25633 : 00000;
25634 : 00000;
25635 : 00000;
25636 : 00000;
25637 : 00000;
25640 : 00000;
25641 : 00000;
25642 : 00000;
25643 : 00000;
25644 : 00000;
25645 : 00000;
25646 : 00000;
25647 : 00000;
25650 : 00000;
25651 : 00000;
25652 : 00000;
25653 : 00000;
25654 : 00000;
25655 : 00000;
25656 : 00000;
25657 : 00000;
25660 : 00000;
25661 : 00000;
25662 : 00000;
25663 : 00000;
25664 : 00000;
25665 : 00000;
25666 : 00000;
25667 : 00000;
25670 : 00000;
25671 : 00000;
25672 : 00000;
25673 : 00000;
25674 : 00000;
25675 : 00000;
25676 : 00000;
25677 : 00000;
25700 : 00000;
25701 : 00000;
25702 : 00000;
25703 : 00000;
25704 : 00000;
25705 : 00000;
25706 : 00000;
25707 : 00000;
25710 : 00000;
25711 : 00000;
25712 : 00000;
25713 : 00000;
25714 : 00000;
25715 : 00000;
25716 : 00000;
25717 : 00000;
25720 : 00000;
25721 : 00000;
25722 : 00000;
25723 : 00000;
25724 : 00000;
25725 : 00000;
25726 : 00000;
25727 : 00000;
25730 : 00000;
25731 : 00000;
25732 : 00000;
25733 : 00000;
25734 : 00000;
25735 : 00000;
25736 : 00000;
25737 : 00000;
25740 : 00000;
25741 : 00000;
25742 : 00000;
25743 : 00000;
25744 : 00000;
25745 : 00000;
25746 : 00000;
25747 : 00000;
25750 : 00000;
25751 : 00000;
25752 : 00000;
25753 : 00000;
25754 : 00000;
25755 : 00000;
25756 : 00000;
25757 : 00000;
25760 : 00000;
25761 : 00000;
25762 : 00000;
25763 : 00000;
25764 : 00000;
25765 : 00000;
25766 : 00000;
25767 : 00000;
25770 : 00000;
25771 : 00000;
25772 : 00000;
25773 : 00000;
25774 : 00000;
25775 : 00000;
25776 : 00000;
25777 : 00000;
END;
